`ifndef END2END_SVH
`define END2END_SVH

//TODO: NEEDS IMPLEMENTATION

`endif