/*
*   Copyright 2016 Purdue University
*   
*   Licensed under the Apache License, Version 2.0 (the "License");
*   you may not use this file except in compliance with the License.
*   You may obtain a copy of the License at
*   
*       http://www.apache.org/licenses/LICENSE-2.0
*   
*   Unless required by applicable law or agreed to in writing, software
*   distributed under the License is distributed on an "AS IS" BASIS,
*   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
*   See the License for the specific language governing permissions and
*   limitations under the License.
*
*
*   Filename:     ooo_decode_stage.sv
*
*   Created by:   Owen Prince
*   Email:        oprince@purdue.edu
*   Date Created: 02/24/2022
*   Description:  Decode stage for out of order pipeline 
*/

`include "ooo_fetch_decode_if.vh"
`include "ooo_decode_execute_if.vh"
`include "control_unit_if.vh"
`include "component_selection_defines.vh"
`include "rv32i_reg_file_if.vh"
`include "ooo_hazard_unit_if.vh"
`include "cache_control_if.vh"
`include "completion_buffer_if.vh"
`include "ooo_bypass_unit_if.vh"

module ooo_decode_stage (
  input logic CLK, nRST, halt, ihit,
  ooo_fetch_decode_if.decode fetch_decode_if,
  ooo_decode_execute_if.decode decode_execute_if,
  rv32i_reg_file_if.decode rf_if,
  ooo_hazard_unit_if.decode hazard_if,
  cache_control_if.pipeline cc_if,
  completion_buffer_if.decode cb_if,
  ooo_bypass_unit_if.decode bypass_if
);

  import rv32i_types_pkg::*;
  import alu_types_pkg::*;
  //import rv32m_pkg::*;
  import machine_mode_types_1_11_pkg::*;

  logic ebreak_ecall;
  logic stall_csr;
  assign ebreak_ecall = cu_if.breakpoint | cu_if.ecall_insn | cu_if.ret_insn;

  // Interface declarations
  control_unit_if   cu_if();
 
  // Module instantiations
  /*******************************************************
  * Input to the Control Unit
  *******************************************************/
  assign cu_if.instr = fetch_decode_if.instr;
  assign decode_execute_if.instr = fetch_decode_if.instr;
  assign cu_if.pc_en = hazard_if.pc_en;
  
  control_unit cu (
    .cu_if(cu_if)
  );
  
  /*******************************************************
  *** fence instruction and Associated Logic 
  *******************************************************/
  // posedge detector for ifence
  // subsequent ifences will have same effect as a single fence
  /*logic ifence_reg;
  logic ifence_pulse;

  always_ff @ (posedge CLK, negedge nRST) begin
    if (~nRST)
      ifence_reg <= 1'b0;
    else if (hazard_if.pc_en)
      ifence_reg <= cu_if.ifence;
  end
  
  assign ifence_pulse = cu_if.ifence && ~ifence_reg;
  assign cc_if.icache_flush = ifence_pulse;
  assign cc_if.icache_clear = 1'b0;
  assign cc_if.dcache_flush = ifence_pulse;
  assign cc_if.dcache_clear = 1'b0; */

  assign hazard_if.ifence_decode = cu_if.ifence;

  //regs to detect flush completion
  /*logic dflushed, iflushed;

  always_ff @ (posedge CLK, negedge nRST) begin
    if (~nRST)
      iflushed <= 1'b1;
    else if (ifence_pulse)
      iflushed <= 1'b0;
    else if (cc_if.iflush_done & hazard_if.pc_en)
      iflushed <= 1'b1;
  end

  always_ff @ (posedge CLK, negedge nRST) begin
    if (~nRST)
      dflushed <= 1'b1;
    else if (ifence_pulse)
      dflushed <= 1'b0;
    else if (cc_if.dflush_done & hazard_if.pc_en)
      dflushed <= 1'b1;
  end
  
  assign hazard_if.dflushed = dflushed;
  assign hazard_if.iflushed = iflushed;
  assign hazard_if.ifence = decode_execute_if.ifence;
  assign hazard_if.ifence_pc = decode_execute_if.pc; */


  /*******************************************************
  * Reg File Logic
  *******************************************************/
  assign rf_if.rs1 = cu_if.reg_rs1;
  assign rf_if.rs2 = cu_if.reg_rs2;

  assign rf_if.rd_decode = cu_if.reg_rd;
  assign rf_if.rden = cu_if.wen & ~cu_if.branch & ~hazard_if.stall_fetch_decode & ~hazard_if.npc_sel & ~stall_csr & ~ebreak_ecall & ~hazard_if.ifence_ex; 
  assign rf_if.clear_status = hazard_if.decode_execute_flush;
  
  /*******************************************************
  *** Sign Extensions of the Immediate Value
  *******************************************************/
  word_t imm_I_ext, imm_S_ext, imm_UJ_ext;

  // for jump calculation
  assign imm_I_ext  = {{20{cu_if.imm_I[11]}}, cu_if.imm_I};
  assign imm_UJ_ext = {{11{cu_if.imm_UJ[20]}}, cu_if.imm_UJ};

  // for source selection
  assign imm_S_ext  = {{20{cu_if.imm_S[11]}}, cu_if.imm_S};
  
  // word_t next_immediate;
  // always_comb begin
    
  // end 



  /*******************************************************
  *** Source Select Logic
  *******************************************************/
  word_t imm_or_shamt, next_reg_file_wdata;
  assign imm_or_shamt = (cu_if.imm_shamt_sel == 1'b1) ? cu_if.shamt : imm_I_ext;

  word_t fu_source_a;
  word_t fu_source_b;
  word_t rs1_data;
  word_t rs2_data;
  assign rs1_data = bypass_if.rs1_bypass_ena ? bypass_if.rs1_bypass_data : rf_if.rs1_data;
  assign rs2_data = bypass_if.rs2_bypass_ena ? bypass_if.rs2_bypass_data : rf_if.rs2_data;
  always_comb begin
    case (cu_if.source_a_sel)
      2'd0: fu_source_a = rs1_data;
      2'd1: fu_source_a = imm_S_ext;
      2'd2: fu_source_a = fetch_decode_if.pc;
      2'd3: fu_source_a = '0; //Not Used 
    endcase
  end
 
  always_comb begin
    case(cu_if.source_b_sel)
      2'd0: fu_source_b = rs1_data;
      2'd1: fu_source_b = rs2_data;
      2'd2: fu_source_b = imm_or_shamt;
      2'd3: fu_source_b = cu_if.imm_U;
    endcase
  end

  always_comb begin
    case(cu_if.arith_sigs.w_src)
      3'd1    : next_reg_file_wdata = fetch_decode_if.pc4;
      3'd2    : next_reg_file_wdata = cu_if.imm_U;
      default : next_reg_file_wdata = '0; 
    endcase
  end
  
  /*******************************************************
  *** Jump Target Calculator and Associated Logic 
  *******************************************************/
  jump_control_signals_t jump_signals;
  word_t base, offset;

  always_comb begin
    if (cu_if.j_sel) begin
      base = fetch_decode_if.pc;
      offset = imm_UJ_ext;
    end else begin
      base = fu_source_a;
      offset = imm_I_ext;
    end
  end 
  assign jump_signals.j_base = base;
  assign jump_signals.j_offset = offset;
  assign jump_signals.jump_instr = cu_if.jump;
  assign jump_signals.j_sel = cu_if.j_sel;
 

  /*******************************************************
  *** Hazard unit connection  
  *******************************************************/
  assign hazard_if.halt = cu_if.halt; //TODO
  assign hazard_if.rs1_busy  = rf_if.rs1_busy & ~bypass_if.rs1_bypass_ena;
  assign hazard_if.rs2_busy  = rf_if.rs2_busy & ~bypass_if.rs2_bypass_ena;
  assign hazard_if.rd_busy   = rf_if.rd_busy;
  assign hazard_if.source_a_sel = cu_if.source_a_sel;
  assign hazard_if.source_b_sel = cu_if.source_b_sel;
  assign hazard_if.fu_type = cu_if.sfu_type;
  always_comb begin
    case (cu_if.sfu_type) 
      LOADSTORE_S: hazard_if.wen = cu_if.lsu_sigs.wen;
      ARITH_S:     hazard_if.wen = cu_if.arith_sigs.wen;
      DIV_S:       hazard_if.wen = cu_if.div_sigs.wen;
      MUL_S:       hazard_if.wen = cu_if.mult_sigs.wen;
    endcase
  end

  /*******************************************************
  *** Bypass Unit logic 
  *******************************************************/
  assign bypass_if.rs1 = cu_if.reg_rs1; 
  assign bypass_if.rs2 = cu_if.reg_rs2; 


  /*********************************************************
  *** Signals for Bind Tracking - Read-Only, These don't affect execution
  *********************************************************/
  // CPU Tracker binding
  cpu_tracker_t CPU_TRACKER;
  assign cb_if.CPU_TRACKER_decode = CPU_TRACKER;
  assign CPU_TRACKER.funct3     = cu_if.instr[14:12];
  assign CPU_TRACKER.funct12    = cu_if.instr[31:20];
  assign CPU_TRACKER.instr_30   = cu_if.instr[30];
  assign CPU_TRACKER.imm_S      = cu_if.imm_S;
  assign CPU_TRACKER.imm_I      = cu_if.imm_I;
  assign CPU_TRACKER.imm_U      = cu_if.imm_U;
  assign CPU_TRACKER.imm_UJ_ext = imm_UJ_ext;
  assign CPU_TRACKER.imm_SB     = cu_if.imm_SB;
  assign CPU_TRACKER.reg_rs1    = cu_if.reg_rs1;
  assign CPU_TRACKER.reg_rs2    = cu_if.reg_rs2;
  assign CPU_TRACKER.instr      = fetch_decode_if.instr;
  assign CPU_TRACKER.reg_rd     = cu_if.reg_rd;
  assign CPU_TRACKER.pc         = fetch_decode_if.pc;
  assign CPU_TRACKER.opcode     = cu_if.opcode;

  /*********************************************************
  *** Stall signals
  *********************************************************/
  assign decode_execute_if.stall_multiply = hazard_if.stall_mu; 
  assign decode_execute_if.stall_divide = hazard_if.stall_du; 
  assign decode_execute_if.stall_arith = hazard_if.stall_au; 
  assign decode_execute_if.stall_loadstore = hazard_if.stall_ls; 

  /*********************************************************
  *** Completion buffer signals
  *********************************************************/
  logic TODO = 0;
  assign cb_if.alloc_ena =  ~hazard_if.stall_fetch_decode && ~hazard_if.npc_sel && cu_if.opcode != MISCMEM & ~ebreak_ecall & ~hazard_if.ifence_ex;
  assign cb_if.rv32v_wb_scalar_ena  = TODO;
  assign cb_if.rv32v_instr  = TODO;
  assign cb_if.opcode = cu_if.opcode;


  /***** CPU_TRACKER, FUNCTIONAL UNIT TYPE LATCH *****/
  always_ff @(posedge CLK, negedge nRST) begin : TOP_CONTROL_SIGNALS
    if (~nRST) begin
      decode_execute_if.sfu_type   <= ARITH_S;
      //decode_execute_if.tracker_sigs <= '0;
    end else begin 
        if ((hazard_if.decode_execute_flush |(hazard_if.stall_fetch_decode & ~hazard_if.stall_ex)) | halt) begin
          decode_execute_if.sfu_type   <= ARITH_S;
          //decode_execute_if.tracker_sigs <= '0;
        end else if(~hazard_if.stall_ex) begin
          decode_execute_if.sfu_type   <= cu_if.sfu_type;
          //decode_execute_if.tracker_sigs <= CPU_TRACKER;
        end
    end
  end


  /***** CSR INSTRUCTION LATCH *****/
  typedef struct packed {
    logic [7:0] vl;
    logic [7:0] vtype;
  } vector_csr_t;

  vector_csr_t vcsr;

  assign vcsr.vtype = cu_if.csr_sigs.vtype_imm ? cu_if.csr_sigs.csr_imm_value[7:0] : rf_if.rs2_data;
  assign vcsr.vl    = cu_if.csr_sigs.vl_imm ? {3'd0, cu_if.reg_rs1} : rf_if.rs1_data[7:0];
  
  assign stall_csr = cu_if.csr_sigs.csr_instr & ~hazard_if.rob_empty & ~hazard_if.csr_flush;
  assign hazard_if.stall_csr = stall_csr;
//  assign decode_execute_if.next_vtype_csr    <= (vcu_if.cfgsel == VSETIVLI) || (vcu_if.cfgsel == VSETVLI) ? {24'd0, vop_c.vma, vop_c.vta, vop_c.sew, vop_c.lmul} : decode_execute_if.xs2;
//  assign decode_execute_if.next_avl_csr      <= (vcu_if.cfgsel == VSETIVLI) ? vcu_if.imm_5 : decode_execute_if.xs1;

  always_ff @(posedge CLK, negedge nRST) begin : CSR_INSTRS
    if (~nRST) begin
      decode_execute_if.csr_sigs <= '0;
    end else begin
      if (hazard_if.decode_execute_flush | stall_csr | hazard_if.csr_ready | (hazard_if.stall_fetch_decode & ~hazard_if.stall_ex)) begin 
        decode_execute_if.csr_sigs <= '0;
      end else if (hazard_if.rob_empty & ~hazard_if.stall_au & ~hazard_if.csr_flush) begin
        // Control signals 
        decode_execute_if.csr_sigs.csr_swap      <= cu_if.csr_sigs.csr_swap;
        decode_execute_if.csr_sigs.csr_clr       <= cu_if.csr_sigs.csr_clr;
        decode_execute_if.csr_sigs.csr_set       <= cu_if.csr_sigs.csr_set;
        decode_execute_if.csr_sigs.csr_addr      <= cu_if.csr_sigs.csr_addr;
        decode_execute_if.csr_sigs.csr_imm       <= cu_if.csr_sigs.csr_imm;
        // Data 
        decode_execute_if.csr_sigs.csr_imm_value <= cu_if.csr_sigs.csr_imm_value;
        decode_execute_if.csr_sigs.csr_instr     <= cu_if.csr_sigs.csr_instr;
        decode_execute_if.csr_sigs.csr_wdata     <= cu_if.csr_sigs.vector_csr_instr ? {8'd0, vcsr} : 
                                                    cu_if.csr_sigs.csr_imm ? cu_if.csr_sigs.csr_imm_value : fu_source_a;
        decode_execute_if.csr_sigs.vector_csr_instr <= cu_if.csr_sigs.vector_csr_instr;
        decode_execute_if.csr_sigs.instr         <= fetch_decode_if.instr;
      end
    end
  end

  /***** HALT INSTRUCTION LATCH *****/
  always_ff @(posedge CLK, negedge nRST) begin : HALT_INSTR
    if (~nRST) begin
            decode_execute_if.halt_instr <= '0;
    end 
    else begin 
        if ((hazard_if.decode_execute_flush |(hazard_if.stall_fetch_decode & ~hazard_if.stall_ex)) | hazard_if.stall_au | hazard_if.stall_mu | hazard_if.stall_du | hazard_if.stall_ls) begin
          decode_execute_if.halt_instr <= '0;
        end else if(~hazard_if.stall_ex & ~(hazard_if.stall_au | hazard_if.stall_mu | hazard_if.stall_du | hazard_if.stall_ls)) begin
          decode_execute_if.halt_instr <= cu_if.halt;
        end
    end
  end

  // Busy signal for decode stage
  assign hazard_if.busy_decode = stall_csr | cu_if.halt & (hazard_if.stall_au | hazard_if.stall_mu | hazard_if.stall_du | hazard_if.stall_ls);

  /***** MULT, DIV, LSU INSTRUCTION LATCH *****/
  always_ff @(posedge CLK, negedge nRST) begin : FUNCTIONAL_UNITS
    if (~nRST) begin
      decode_execute_if.mult_sigs <= '0;
      decode_execute_if.div_sigs <= '0;
      decode_execute_if.lsu_sigs <= '0;
    end else begin
      if (hazard_if.decode_execute_flush | (hazard_if.stall_fetch_decode & ~hazard_if.stall_ex) | halt) begin : FLUSH
        decode_execute_if.mult_sigs <= '0;
        decode_execute_if.div_sigs <= '0;
        decode_execute_if.lsu_sigs <= '0;
      end else begin
        //MULTIPLY
        if(~cu_if.mult_sigs.ena) begin
          decode_execute_if.mult_sigs <= '0;
        end else if(~(hazard_if.stall_mu) & ~hazard_if.stall_ex) begin
          decode_execute_if.mult_sigs.ena <= cu_if.mult_sigs.ena;
          decode_execute_if.mult_sigs.high_low_sel <= cu_if.mult_sigs.high_low_sel;
          decode_execute_if.mult_sigs.is_signed <= cu_if.mult_sigs.is_signed;
          decode_execute_if.mult_sigs.decode_done <= cu_if.mult_sigs.decode_done;
          decode_execute_if.mult_sigs.wen <= cu_if.mult_sigs.wen;
          decode_execute_if.mult_sigs.reg_rd <= cu_if.mult_sigs.reg_rd;
          decode_execute_if.mult_sigs.ready_mu <= cu_if.mult_sigs.ready_mu;
          decode_execute_if.mult_sigs.index_mu <= cb_if.cur_tail;
        end
       
        //DIVIDE
        if(~cu_if.div_sigs.ena) begin
          decode_execute_if.div_sigs <= '0;
        end else if(~(hazard_if.stall_du) & ~hazard_if.stall_ex) begin
        //if(~(hazard_if.stall_du)) begin
          decode_execute_if.div_sigs.ena <= cu_if.div_sigs.ena;
          decode_execute_if.div_sigs.div_type <= cu_if.div_sigs.div_type;
          decode_execute_if.div_sigs.is_signed <= cu_if.div_sigs.is_signed;
          decode_execute_if.div_sigs.wen <= cu_if.div_sigs.wen;
          decode_execute_if.div_sigs.reg_rd <= cu_if.div_sigs.reg_rd;
          decode_execute_if.div_sigs.ready_du <= cu_if.div_sigs.ready_du;
          decode_execute_if.div_sigs.index_du <= cb_if.cur_tail;
        end

        // LOADSTORE
        if(~cu_if.lsu_sigs.ena) begin
          decode_execute_if.lsu_sigs <= '0;
        end else if(~(hazard_if.stall_ls) & ~hazard_if.stall_ex) begin
          decode_execute_if.lsu_sigs.load_type <= cu_if.lsu_sigs.load_type;
          //decode_execute_if.lsu_sigs.byte_en <= cu_if.lsu_sigs.byte_en;
          decode_execute_if.lsu_sigs.dren <= cu_if.lsu_sigs.dren;
          decode_execute_if.lsu_sigs.dwen <= cu_if.lsu_sigs.dwen;
          decode_execute_if.lsu_sigs.opcode <= cu_if.lsu_sigs.opcode;
          decode_execute_if.lsu_sigs.wen <= cu_if.lsu_sigs.wen;
          decode_execute_if.lsu_sigs.reg_rd <= cu_if.lsu_sigs.reg_rd;
          decode_execute_if.lsu_sigs.ready_ls <= cu_if.lsu_sigs.ready_ls;
          decode_execute_if.lsu_sigs.index_ls <= cb_if.cur_tail;
          decode_execute_if.store_data <= rs2_data;
        end

      end
    end
  end

  /***** FUNCTIONAL UNIT SOURCE LATCHES *****/
  always_ff @(posedge CLK, negedge nRST) begin : SOURCE_LATCHES
    if(~nRST) begin
      decode_execute_if.pc <= '0;
      decode_execute_if.pc4 <= '0;
      decode_execute_if.immediate <= '0;
      decode_execute_if.port_a <= '0; 
      decode_execute_if.port_b <= '0; 
      decode_execute_if.lsu_sigs.opcode <= '0;    
      decode_execute_if.ifence <= '0;    
    end else begin 
      if(hazard_if.decode_execute_flush | (hazard_if.stall_fetch_decode & ~hazard_if.stall_ex) | halt) begin
        decode_execute_if.pc <= '0;
        decode_execute_if.pc4 <= '0;
        decode_execute_if.immediate <= '0;
        decode_execute_if.port_a <= '0; 
        decode_execute_if.port_b <= '0; 
        decode_execute_if.lsu_sigs.opcode <= '0;
        decode_execute_if.ifence <= '0;    
      end else if(~hazard_if.stall_ex) begin
        decode_execute_if.pc <= fetch_decode_if.pc;
        decode_execute_if.pc4 <= fetch_decode_if.pc4;
        decode_execute_if.immediate <= cu_if.imm_SB; // TODO figure out how to do this
        decode_execute_if.port_a <= fu_source_a; 
        decode_execute_if.port_b <= fu_source_b; 
        decode_execute_if.lsu_sigs.opcode <= cu_if.opcode;
        decode_execute_if.ifence <= cu_if.ifence;    
      end
    end
  end

  /***** ARITHMETIC UNIT/CSR/EXCEPTION LATCH *****/
  always_ff @(posedge CLK, negedge nRST) begin : ARITH_UNIT
    if (~nRST) begin
      decode_execute_if.arith_sigs <= '0;
      decode_execute_if.reg_file_wdata <= '0;
      //JUMP
      decode_execute_if.jump_sigs        <= '0;
      //BRANCH
      decode_execute_if.branch_sigs <= '0;
      //Exceptions
      decode_execute_if.exception_sigs <= '0;
        
    end else begin
      if (hazard_if.decode_execute_flush | (~hazard_if.stall_ex & hazard_if.stall_fetch_decode) | halt) begin
        decode_execute_if.arith_sigs <= '0;
        decode_execute_if.reg_file_wdata <= '0;
        //JUMP
        decode_execute_if.jump_sigs <= '0;
        //BRANCH
        decode_execute_if.branch_sigs <= '0;
        //Exceptions
        decode_execute_if.exception_sigs <= '0;

      end else if(~cu_if.arith_sigs.ena & ~hazard_if.stall_ex) begin
        decode_execute_if.arith_sigs <= '0;
        decode_execute_if.reg_file_wdata <= next_reg_file_wdata;
        decode_execute_if.jump_sigs <= '0;
        decode_execute_if.branch_sigs <= 0;

        //Exceptions
        // elaborateed because half of the signals are form cu_if and 
        // other half is from the fetch decode latch
        decode_execute_if.exception_sigs.illegal_insn <= cu_if.illegal_insn;
        decode_execute_if.exception_sigs.breakpoint   <= cu_if.breakpoint;
        decode_execute_if.exception_sigs.ecall_insn   <= cu_if.ecall_insn;
        decode_execute_if.exception_sigs.ret_insn     <= cu_if.ret_insn;
        decode_execute_if.exception_sigs.token        <= fetch_decode_if.token;
        decode_execute_if.exception_sigs.mal_insn     <= fetch_decode_if.mal_insn;
        decode_execute_if.exception_sigs.fault_insn   <= fetch_decode_if.fault_insn;
        decode_execute_if.exception_sigs.wfi          <= cu_if.wfi;
        decode_execute_if.exception_sigs.w_src        <= cu_if.arith_sigs.w_src;
      end else if(~hazard_if.stall_au & ~hazard_if.stall_ex) begin
        decode_execute_if.arith_sigs.ena <= cu_if.arith_sigs.ena;
        decode_execute_if.arith_sigs.alu_op <= cu_if.arith_sigs.alu_op;
        decode_execute_if.arith_sigs.w_src <= cu_if.arith_sigs.w_src;
        decode_execute_if.arith_sigs.wen <= cu_if.arith_sigs.wen;
        decode_execute_if.arith_sigs.reg_rd <= cu_if.arith_sigs.reg_rd;
        decode_execute_if.arith_sigs.ready_a <= cu_if.arith_sigs.ready_a;
        decode_execute_if.arith_sigs.index_a <= cb_if.cur_tail;

        decode_execute_if.reg_file_wdata <= next_reg_file_wdata;
        //JUMP
        decode_execute_if.jump_sigs <= jump_signals;
        //BRANCH
        // pretty sure this line is unecessary
        // decode_execute_if.branch_sigs.br_imm_sb       <= cu_if.imm_SB;
        decode_execute_if.branch_sigs.branch_type  <= cu_if.branch_type;
        decode_execute_if.branch_sigs.branch_instr      <= cu_if.branch;
        //BRANCH PREDICTOR UPDATE
        decode_execute_if.branch_sigs.prediction <= fetch_decode_if.prediction;

        //Exceptions
        // elaborateed because half of the signals are form cu_if and 
        // other half is from the fetch decode latch
        decode_execute_if.exception_sigs.illegal_insn <= cu_if.illegal_insn;
        decode_execute_if.exception_sigs.breakpoint   <= cu_if.breakpoint;
        decode_execute_if.exception_sigs.ecall_insn   <= cu_if.ecall_insn;
        decode_execute_if.exception_sigs.ret_insn     <= cu_if.ret_insn;
        decode_execute_if.exception_sigs.token        <= fetch_decode_if.token;
        decode_execute_if.exception_sigs.mal_insn     <= fetch_decode_if.mal_insn;
        decode_execute_if.exception_sigs.fault_insn   <= fetch_decode_if.fault_insn;
        decode_execute_if.exception_sigs.wfi          <= cu_if.wfi;
        decode_execute_if.exception_sigs.w_src        <= cu_if.arith_sigs.w_src;

      end
    end
  end

  //assign hazard_if.instr_wait_ihit = cu_if.branch | cu_if.jump | cu_if.csr_sigs.csr_instr;
  //assign hazard_if.instr_wait_ihit = 1;

  logic [18:0] write_conflict_reg, next_write_conflict_reg;
  logic div_write_conflict_stall;
  logic mul_write_conflict_stall;
  logic alu_write_conflict_stall;
  logic write_conflict_stall;
  logic div_special_case;
  logic alu_ena;

  assign hazard_if.wb_port_conflict  = write_conflict_stall;

  assign alu_ena = cu_if.arith_sigs.ena | cu_if.illegal_insn | fetch_decode_if.mal_insn;
  assign div_write_conflict_stall = cu_if.div_sigs.ena & div_special_case ? write_conflict_reg[0] :
                                    cu_if.div_sigs.ena ? write_conflict_reg[17] :
                                    0;
  assign mul_write_conflict_stall = cu_if.mult_sigs.ena & write_conflict_reg[3];
  assign alu_write_conflict_stall = cu_if.csr_sigs.csr_instr ? write_conflict_reg[1] :
                                    alu_ena ? write_conflict_reg[0] :
                                    0;
  assign write_conflict_stall     = (div_write_conflict_stall | mul_write_conflict_stall | alu_write_conflict_stall) & ~ebreak_ecall & (cu_if.opcode != opcode_t'('h0));
  assign div_special_case         = fu_source_a == 32'h8000_0000 | fu_source_b == 32'hffff_ffff | fu_source_b == 32'h0;       

  always_ff @(posedge CLK, negedge nRST) begin
    if (~nRST) begin
        write_conflict_reg <= '0;
    end else if (~hazard_if.stall_fetch_decode) begin
        write_conflict_reg <= next_write_conflict_reg >> 1;
    end else begin
        write_conflict_reg <= write_conflict_reg >> 1;
    end
  end

  always_comb begin
    next_write_conflict_reg = write_conflict_reg;
    if (cu_if.div_sigs.ena) begin
        if (div_special_case) next_write_conflict_reg = write_conflict_reg | 1'b1;
        else next_write_conflict_reg = write_conflict_reg | 18'b100000000000000000;
    end else if (cu_if.mult_sigs.ena) begin
        next_write_conflict_reg = write_conflict_reg | 4'b1000;
    end else if (cu_if.csr_sigs.csr_instr) begin
        next_write_conflict_reg = write_conflict_reg | 2'b10;
    end else if (alu_ena) begin
        next_write_conflict_reg = write_conflict_reg | 1'b1;
    end
  end

endmodule
