`ifndef DUT_PARAMS_SVH
`define DUT_PARAMS_SVH

package dut_params;

localparam NUM_CPUS_USED 2;
localparam BLOCK_SIZE_WORDS 2;
localparam WORD_W 32;

endpackage
`endif
