`timescale 1ns/100ps
module tb_FPU_top_level();
   reg clk = 0;
   reg nrst;
   reg [31:0] floating_point1;
   reg [31:0] floating_point2;
   reg [2:0]  frm;
   reg [31:0] floating_point_out;
   reg [6:0]  funct7;
   reg [4:0]  flags;
   
   always begin
      clk = ~clk;
      #1;
   end

   FPU_top_level DUT (
		      .clk(clk),
		      .nrst(nrst),
		      .floating_point1(floating_point1),
		      .floating_point2(floating_point2),
		      .frm(frm),
		      .funct7(funct7),
		      .floating_point_out(floating_point_out),
		      .flags(flags)
		      );
   
   shortreal        result_real;
   reg  [31:0] result_binary;
   shortreal        fp1_real;
   shortreal        fp2_real;
   shortreal        fp_out_real;
   shortreal        fp_exp;
   shortreal        fp_frac;
   int       i;
   int       j = 0;
   //real val1;
   //shortreal val2;
   
   task random_check;
      begin
         //$display($bits(val1));
   	 //$display($bits(val2));
  //subnormal number
	 frm = $random() % 8;
	 //frm       = 3'b000;
	 //frm = 3'b111;
	 //funct7 = 7'b0100000;
	 funct7 = 7'b0100100;
	 floating_point1 = $random(); //0
	 floating_point2 = $random(); //10010001110111111110100000100011
	 //Error: expected = 0 00011101 00110010000000000000000, 
         //	calculated = 0 00100001 00010011001000000000000,
	 /*if (i == 0) begin
	 floating_point1 = 32'b01000001000111000000000000000000; //9.75
	 floating_point2 = 32'b00111111000100000000000000000000; //0.5625
	 //Error: expected = 0 10000010  00100110000000000000000, 
	 //	calculated = 0 10000010 10010011000000000000000
	 end else if (i == 1) begin
         floating_point1 = 32'b01000010101110010110011001100110; //92.7
	 floating_point2 = 32'b01000001110110110011001100110011; //27.4
	 //Error: expected = 0 10000101  00000101001100110011001, 
	 //	calculated = 0 10000101 10000010100110011001100
	 end else if (i == 2) begin
	 floating_point1 = 32'b01000101100011110101110101100010; //4587.673
         floating_point2 = 32'b01000011111100111101011000101011; //487.6732
	 //Error: expected = 0 10001011  00000000001111111111111, 
	 //	calculated = 0 10001011 10000000000111111111111
	 end else if (i == 3) begin
	 floating_point1 = 32'b01001011000100110011000110001111; //9646479.12357
         floating_point2 = 32'b01000111111100010010011111010110; //123471.6732
	 end else if (i == 4) begin
	 floating_point1 = 32'b01000111001101101011010001101010; //46772.414
         floating_point2 = 32'b01000101000100111111011001100110; //2367.4
	 end else if (i == 5) begin
         floating_point1 = 32'b11000001000111000000000000000000; //-9.75
	 floating_point2 = 32'b10111111000100000000000000000000; //-0.5625
	 //Error: expected = 11000001000100110000000000000000, 
	 //	calculated = 11000001000100101111111111111111,     1+

	 //Error: expected = 1 10000010 00100110000000000000000, 
	 //	calculated = 1 10000011  01101101000000000000000,
	 end else if (i == 6) begin
         floating_point1 = 32'b11000010101110010110011001100110; //-92.7
	 floating_point2 = 32'b11000001110110110011001100110011; //-27.4
	 end else if (i == 7) begin
	 floating_point1 = 32'b11000101100011110101110101100010; //-4587.673
         floating_point2 = 32'b11000011111100111101011000101011; //-487.6732
	 end else if (i == 8) begin
	 floating_point1 = 32'b11001011000100110011000110001111; //-9646479.12357
         floating_point2 = 32'b11000111111100010010011111010110; //-123471.6732
	 end else if (i == 9) begin
	 floating_point1 = 32'b11000111001101101011010001101010; //-46772.414
         floating_point2 = 32'b11000101000100111111011001100110; //-2367.4
	 end else if (i == 10) begin
	 floating_point1 = 32'b00111111000100000000000000000000; //0.5625
         floating_point2 = 32'b01000001000111000000000000000000; //9.75
	 end else if (i == 11) begin
	 floating_point1 = 32'b01000001110110110011001100110011; //27.4
         floating_point2 = 32'b01000010101110010110011001100110; //92.7
	 end else if (i == 12) begin
         floating_point1 = 32'b01000011111100111101011000101011; //487.6732
	 floating_point2 = 32'b01000101100011110101110101100010; //4587.673
	 end else if (i == 13) begin
         floating_point1 = 32'b01000111111100010010011111010110; //123471.6732
	 floating_point2 = 32'b01001011000100110011000110001111; //9646479.12357
	 end else if (i == 14) begin
         floating_point1 = 32'b01000101000100111111011001100110; //2367.4
	 floating_point2 = 32'b01000111001101101011010001101010; //46772.414
	 end else if (i == 15) begin
	 floating_point1 = 32'b00111110100000000000000000000000; //.25
	 floating_point2 = 32'b01000010110010000000000000000000; //100
	 end else if (i == 16) begin
	 floating_point1 = 32'b11000001110110110011001100110011; //-27.4
         floating_point2 = 32'b11000010101110010110011001100110; //-92.7
	 end else if (i == 17) begin
	 floating_point1 = 32'b11000101000100100011011001100110; //-2367.3999
	 floating_point2 = 32'b11000111001110101011010101101010; //-46773.4141
	 end else if (i == 18) begin
         floating_point1 = 32'b11000010100100011111111101111101; //-72.999
	 floating_point2 = 32'b11001110001100100110011001001001; //-748261946.14893
	 end else if (i == 19) begin
	 floating_point1 = 32'b11000010110101101101011100001010; //-107.42
	 floating_point2 = 32'b11000111101110111110011110001110; //-96207.111
	 end else if (i == 20) begin
	 floating_point1 = 32'b10111111000100000000000000000000; //-0.5625
         floating_point2 = 32'b11000001000111000000000000000000; //-9.75
	 //Error: expected = 01000001000100110000000000000000, 
	 //	calculated = 01000001000100101111111111111111 1+
	 end /*else if (i == 21) begin
	 floating_point1 = 32'b01111111100000000000000000000000; //Inf
	 floating_point2 = 32'b11000010101010000011011111001111; //-94.109
 	 end else if (i == 22) begin
         floating_point1 = 32'b11111111100000000000000000000000; //-Inf
	 floating_point2 = 32'b11000001000001101001001100001100; //-8.4109
	 end else if (i == 23) begin
	 floating_point1 = 32'b11000010101010000011011111001111; //-94.109
	 floating_point2 = 32'b01111111100000000000000000000000; //Inf
 	 end else if (i == 24) begin
         floating_point1 = 32'b11000001000001101001001100001100; //-8.4109
	 floating_point2 = 32'b11111111100000000000000000000000; //-Inf
	 end*/ /*else if (i == 25) begin
	 floating_point1 = 32'b11000010101010000011011111001111; //-94.109
	 floating_point2 = 32'b10000000000000000000000000000000; //-0
 	 end else if (i == 26) begin
         floating_point1 = 32'b11000010101010000011011111001111; //-94.109
	 floating_point2 = 32'b00000000000000000000000000000000; //0
	 end else if (i == 27) begin
	 floating_point1 = 32'b11111111100000000000000000000000; //-Inf
	 floating_point2 = 32'b10000000000000000000000000000000; //-0
 	 end else if (i == 28) begin
	 floating_point1 = 32'b10000000000000000000000000000000; //-0
	 floating_point2 = 32'b11000010101110010110011001100110; //-92.7
 	 end else if (i == 29) begin
	 floating_point1 = 32'b00000000000000000000000000000000; //0
	 floating_point2 = 32'b11000010101110010110011001100110; //-92.7
	 end else if (i == 30) begin
         floating_point1 = 32'b11000000100010010101111010000001; //-4.29
	 floating_point2 = 32'b10000100100001001101011000001001; //-3.13e-36
	 end else if (i == 31) begin
         floating_point1 = 32'b01100000101100010111010111000001; //1.023e20
	 floating_point2 = 32'b11100010111001010111010011000101; //-2.11636e21
         end else if (i == 32) begin
         floating_point1 = 32'b01010101011110000100010110101010; //1.71e13
	 floating_point2 = 32'b11001110110011001100110010011101; //-1717980800
	 end else if (i == 33) begin
         floating_point1 = 32'b01100011010010111111100111000110; //3.763e21
	 floating_point2 = 32'b01010111000101010001001110101110; //1.639e14
	 end else if (i == 34) begin
         floating_point1 = 32'b00110101100111111101110101101011; //1.19e-6
	 floating_point2 = 32'b11101010101001100010101011010101; //-1.0044e26
 	 end else if (i == 35) begin
         floating_point1 = 32'b00000101011100111000011100001010; //1.145e-35
	 floating_point2 = 32'b11000000001110110010001010000000; //-2.924
	 end else if (i == 36) begin
         floating_point1 = 32'b00100000110001001011001101000001; //3.332e-19
	 floating_point2 = 32'b11101100010010110011010011011000; //-9.83e26
	 end else if (i == 37) begin
         floating_point1 = 32'b10001101001001001111011000011010; //-5.08e-31
	 floating_point2 = 32'b11011100111100000000000010111001; //-5.4e17 
	 end else if (i == 38) begin
         floating_point1 = 32'b10011100011011011110011000111000; //-7.87e-22
	 floating_point2 = 32'b10111100110011111010100001111001; //-0.0253488887101 
	 //Error: expected = 00111100110011111010100001111001, 
	 //	calculated = 00111100110011111010100001111000   1+
 	 end else if (i == 39) begin
         floating_point1 = 32'b10111010101100010100100001110101; //-0.00135256221984
	 floating_point2 = 32'b11000111111010000101011010001111; //-118957.117188
	 end else if (i == 40) begin
         floating_point1 = 32'b10110110101001000010011001101101; //-4.89e-6
	 floating_point2 = 32'b10111011010001011110001001110110; //-0.00302 
	 end else if (i == 41) begin
         floating_point1 = 32'b11001101010111101011110010011010; //-233556384
	 floating_point2 = 32'b11111110110111110111001011111101; //-1.485e38 
	 end else if (i == 42) begin
         floating_point1 = 32'b10010111100110011010100000101111; //-9.93e-25
	 floating_point2 = 32'b11011001110100101001001010110011; //-7.41e15 //
	 //Error: expected = 01011001110100101001001010110011, 
	 //	calculated = 01011001110100101001001010110010,   1+
	 end else if (i == 43) begin
         floating_point1 = 32'b10010110100100000000010000101101; //-2.3267e-25
	 floating_point2 = 32'b11100011110001010011000011000111; //-7.275e21 //
	 end else if (i == 44) begin
         floating_point1 = 32'b11001111011000111101101010011110; //-3822755328.0
	 floating_point2 = 32'b11111110111100000110010011111101; //-1.5977e+38 //
	 end else if (i == 45) begin
         floating_point1 = 32'b10111000010101011100010001110000; //-5.0966e-5
	 floating_point2 = 32'b10111001111101010000010001110011; //-0.000467333564302
	 //Error: expected = 00111001110110100100101111100101, 
	 //	calculated = 00111001110110100100101111100100   1+
	 end else if (i == 46) begin
         floating_point1 = 32'b10001001001101110101001000010010; //-2.21e-33
	 floating_point2 = 32'b00000000111100111110001100000001; //2.24e-38 
	 end else if (i == 47) begin
         floating_point1 = 32'b10011110001100010100110000111100; //-9.386e-21
	 floating_point2 = 32'b01111001011010001011110111110010; //7.553e34 
	 //Error: expected = 1 11110010 11010001011110111110010, 
	 //	calculated = 1 11110010 00101110100001000001101   neg
	 //		     1 11110010 00101110100001000001110
	 //		     1 11110010 00101110100001000001110
	 end else if (i == 48) begin
         floating_point1 = 32'b11000100100010100001001010001001; //-1104.579
	 floating_point2 = 32'b01110101110001010000110111101011; //4.996e32
	 //Error: expected = 1 11101011 10001010000110111101011, 
 	 //	calculated = 1 11101011 01110101111001000010100   neg
	 end else if (i == 49) begin 
         floating_point1 = 32'b11110001101100110100110011100011;   //-1.77570454712e+30 ssd
	 floating_point2 = 32'b11110010100110011110110011100101;   //-6.09761208551e+30
	 //Error: expected = 0 11100100  10110100011001101011000, 
	 //	calculated = 0 11100101 11011010001100110101100   1e+1s
	 end else if (i == 50) begin 
         floating_point1 = 32'b11110001001101111111001011100010;   //-9.10870145608e+29 ssd
	 floating_point2 = 32'b11110001100111000111000011100011;   //-1.54931626244e+30
	 //Error: expected = 0 11100010  00000001110111011100100, 
	 //	calculated = 0 11100011 10000000111011101110010   1e+1s
	 end else if (i == 51) begin 
         floating_point1 = 32'b11001010000011100100010010010100;   //-2330917.0 ssd
	 floating_point2 = 32'b11001001011000011110010010010010;   //-925257.125
	 //Error: expected = 1 10010011  01010111001011011011111, 
	 //	calculated = 1 10010100 10101011100101101110000   1e+1s
	 end else if (i == 52) begin 
         floating_point1 = 32'b10100110011000110110001001001100;  //-7.88896629161e-16 ssd
	 floating_point2 = 32'b10101001100000011001010001010011;  //-5.7544809575e-14
	 //Error: expected = 0 01010010  11111111001101100011100, 
	 //	calculated = 0 01010011 11111111100110110001110   1e+1s
	 end else if (i == 53) begin 
         floating_point1 = 32'b11100100100000100100110011001001;  //-1.92288774656e+22 ssd
	 floating_point2 = 32'b11100100110110000010000011001001;  //-3.18948731152e+22
	 //Error: expected = 0 11001000  01010111010100000000000, 
	 //	calculated = 0 11000111 10101110101000000000000   1e+1s
	 end else if (i == 54) begin 
         floating_point1 = 32'b10110110001011011000010001101100;  //-2.58560885413e-06 ssd
	 floating_point2 = 32'b10110101110001011100000001101011;  //-1.47336447753e-06
	 //Error: expected = 1 01101011  00101010100100001101101, 
	 //	calculated = 1 01101100 10010101010010000110111   1e+1s
	 end else if (i == 55) begin 
 	 floating_point1 = 32'b11010001010010001000111010100010;  // -53836652544.0 ssd
	 floating_point2 = 32'b11010011000001011101100010100110;  // -5.74865408e+11
	 //Error: expected = 0 10100101  11100101001111101110111, 
	 //	calculated = 0 10100110 11110010100111110111011   1e+1s
	 end else if (i == 56) begin
         floating_point1 = 32'b01100001100111110010000111000011;  //3.66933136993e+20
	 floating_point2 = 32'b01100000100000000111011111000001;  //7.40566381186e+19
	 //Error: expected = 0 11000010  11111100000011110100101, 
	 //	calculated = 0 11000011 11111110000001111010010   1e+1s
	 end else if (i == 57) begin
         floating_point1 = 32'b01010010101011010101001110100101;  //3.72216332288e+11
	 floating_point2 = 32'b01010010010010001100100110100100;  //2.1559410688e+11
	 //Error: expected = 0 10100100  00100011101110110100110, 
	 //	calculated = 0 10100101 10010001110111011010011   1e+1s
	 end else if (i == 58) begin
         floating_point1 = 32'b00101010001011111111010101010100;  //1.56282376363e-13
	 floating_point2 = 32'b00101010010101100101111101010100;  //1.90400917689e-13
	 end else if (i == 59) begin
         floating_point1 = 32'b10101000101110110000110001010001;  //-2.07665119503e-14
	 floating_point2 = 32'b10101000111000011110111001010001;  //-2.50833713202e-14
	 //Error: expected = 0 01001111 00110111000100000000000, 
	 //	calculated = 0 01001111 00110111000011111111111   1+
	 end else if (i == 60) begin
         floating_point1 = 32'b01010101011110011011011110101010;  //1.71604516536e+13
	 floating_point2 = 32'b01010101010100111011000110101010;  //1.45475009249e+13
	 end else if (i == 61) begin
         floating_point1 = 32'b00001001100011100010110100010011;  //3.42276441045e-33
	 floating_point2 = 32'b00001001110010000011010100010011;  //4.81981593651e-33	
	 //Error: expected = 1 0001000111010000010000000000000, 
	 //	calculated = 1 0001000111010000001111111111111 1+
	 end else if (i == 62) begin
         floating_point1 = 32'b10100111001011000000111001001110;  //-2.38775496161e-15 ssd
	 floating_point2 = 32'b00101000011000100100101101010000;  //1.25618509735e-14
	 //Error: expected = 1 01010001 00001101010011101110001, 
	 //	calculated = 1 01010000 11100101011000100011101

	 //Error: expected = 1 01010001 00001101010011101110001, 
	 //	calculated = 1 01010000  11100101011000100011101
	 //			         00011010100111011100010
	 end//*/


         /*
	Error: expected = 1 0010110 010110110111101100101011, /1
	     calculated = 1 0010110 010110110111101100101101, 
	fp1 is = 00000011110101100010011100000111,  1.25867497925e-36
	fp2 is = 00010110010110110111101100101100,  1.77295453068e-25

	Error: expected = 0 11111100 01001001001000111111011, /2
	     calculated = 0 11111100 01001001001000111111101,  
	fp1 is = 01111110001001001001000111111100, 
	fp2 is = 01101110000111100001111111011100,

	Error: expected = 0 11010100 01011000001001111010011, /3
	     calculated = 0 11010100 01011000001001111010101,
	fp1 is = 01101010001011000001001111010100, 
	fp2 is = 01010010001110010111110110100100, 

	Error: expected = 1 01001100 11001100001000101001011,
	     calculated = 1 01001100 11001100001000101001101 /19
	fp1 is = 00010000101011101110101100100001, 
	fp2 is = 00100110011001100001000101001100,

	Error: expected = 1 01001110 01000000110001101001101, /4
	     calculated = 1 01001110 01000000110001101001111, 
	fp1 is = 00010111101111011000011100101111, 
	fp2 is = 00100111001000000110001101001110,

	Error: expected = 0 11110100 11010101111010111110011, 
	     calculated = 0 11110100 11010101111010111110101,  /8
	fp1 is = 01111010011010101111010111110100,
	fp2 is = 01101000000101011101100111010000,

	Error: expected = 0 01010010 10011000010101101010001, 
	     calculated = 0 01010010 10011000010101101010011, /9
	fp1 is = 00101001010011000010101101010010, 
	fp2 is = 00011010000011101100011100110100, 

	Error: expected = 0 01010111 01001101011000101010110, 
	     calculated = 0 01010111 01001101011000101011000, /10
	fp1 is = 00101011101001101011000101010111, 
	fp2 is = 00011001110011111110101100110011,

	Error: expected = 1 11000110 11010100100001111000101,
	     calculated = 1 11000110 11010100100001111000111, /14
	fp1 is = 01001000101101000000100110010001,
	fp2 is = 01100011011010100100001111000110,

	Error: expected = 0 01000011 00000001011000101000010, 
	     calculated = 0 01000011 00000001011000101000100, /17 
	fp1 is = 00100001100000001011000101000011,
	fp2 is = 00001100001110001110101100011000, 

	Error: expected = 0 11001000 01010111010100000000000,  
	     calculated = 0 11000111  10101110101000000000000,  
	fp1 is = 11100100100000100100110011001001,  -1.92288774656e+22
	fp2 is = 11100100110110000010000011001001,  -3.18948731152e+22		//4 329 ss?
Error: expected =  0 11001000 01010111010100000000000, 
     calculated =  0 11001010 01010111010100000000000 
//10w 67

	Error: expected = 0 01001111  00110111000100000000000, 
	     calculated = 0 01010000 10011011100010000000000, 
	fp1 is = 10101000101110110000110001010001,-2.07665119503e-14
	fp2 is = 10101000111000011110111001010001 -2.50833713202e-14

	Error: expected = 1 10010011  01010111001011011011111, 
	     calculated = 1 10010100 10101011100101101101111,  
	fp1 is = 11001010000011100100010010010100, 	-2330917.0
	fp2 is = 11001001011000011110010010010010, 	-925257.125	///1 375

	Error: expected = 1 01101011 00101010100100001101101,
	     calculated = 1 01101100 10010101010010000110110, 
			  1 01101011 00101010100100001101100
	fp1 is = 10110110001011011000010001101100, 	-2.58560885413e-06
	fp2 is = 10110101110001011100000001101011, 	-1.47336447753e-06	///2 396

	Error: expected = 0 10100100  00100011101110110100110,
	     calculated = 0 10100101 10010001110111011010011    
	fp1 is = 01010010101011010101001110100101,	3.72216332288e+11
	fp2 is = 01010010010010001100100110100100,	2.1559410688e+11 ///4 762

	Error: expected = 0 01010010  11111111001101100011100,
	     calculated = 0 01010011 11111111100110110001110, 
	fp1 is = 10100110011000110110001001001100, 	   -7.88896629161e-16
	fp2 is = 10101001100000011001010001010011,	   -5.7544809575e-14   ///5 847
				    1111111110011011000111010

	Error: expected = 0 11000010  11111100000011110100101, 
	     calculated = 0 11000011 11111110000001111010011 
	fp1 is = 01100001100111110010000111000011, 	3.66933136993e+20
	fp2 is = 01100000100000000111011111000001,	7.40566381186e+19      ///6 861

	Error: expected = 0 10100101  11100101001111101110111, 
	     calculated = 0 10100110 11110010100111110111100, 
	fp1 is = 11010001010010001000111010100010, 	53836652544
	fp2 is = 11010011000001011101100010100110	-5.74865408e+11      ///7 1049

	Error: expected = 0 11100010  00000001110111011100100,
	     calculated = 0 11100011 10000000111011101110010,
	 		  0 11100010  00000001110111011100011
	fp1 is = 11110001001101111111001011100010, 	-9.10870145608e+29
	fp2 is = 11110001100111000111000011100011,	-1.54931626244e+30	      ///8 1067

	Error: expected = 0 11100100  10110100011001101011000,
	     calculated = 0 11100101 11011010001100110101100 
	fp1 is = 11110001101100110100110011100011, 	-1.77570454712e+30
	fp2 is = 11110010100110011110110011100101, 	-6.09761208551e+30      ///9 1175

	Error: expected = 0 00100000  10010110010011100100010, 
	     calculated = 0 00100001 11001011001001110010001	///10 1255
	fp1 is = 00010000110100000000101100100001, 
	fp2 is = 00010000010101001110111100100000

	Error: expected = 1 10010100  11010010101001010010110, 
	     calculated = 1 10010101 11101001010100101001011   ///11 1348
	fp1 is = 11001010111100011111111010010101, 
	fp2 is = 11001010011110101010101010010100

	Error: expected = 1 11110111  10111100011101111110010, 
	     calculated = 1 11111000 11011110001110111111001   ///12 1461
	fp1 is = 01111010100001110111111111110101, 
	fp2 is = 01111100000000000000110111111000

	Error: expected = 1 00001111  11010100010110000011001,  ///14 1685
	     calculated = 1 00010000 11101010001011000001101

	Error: expected = 1 01011011    10101111110010101111100,  /////13 1628
	     calculated = 1 01011110 00110101111110010101111
	fp1 is = 00101110111001101110100101011101, 
	fp2 is = 00101111000011100111000101011110

	Error: expected = 0 11001111 11010011101000000011011, 
	     calculated = 0 11001111 11010011101000000011101   /// 1908
	fp1 is = 0 11001111 11010011100110111001111,  2.20821577793e+24
	fp2 is = 1 11000001 00100110011011011000001   -8.48630254245e+19

	Error: expected = 0 10111011 01001010110101010111011, 
	     calculated = 0 10111011 01001010110101010111101  /// 2192
	fp1 is = 0 10100011 10011011110100110100011, 
	fp2 is = 1 10111011 01001010110101010111011


	Error: expected = 1 01011011    10101111110010101111100, 
	     calculated = 1 01011110 00110101111110010101111   // 1628
			  1 01011011 01101011111100101011110
	fp1 is = 0 01011101 11001101110100101011101,  1.05006427165e-10
	fp2 is = 0 01011110 00011100111000101011110   1.2955100881e-10


	Error: expected = 0 11101001   01001101111100111011000, 
	     calculated = 0 11101011 01010011011111001110110  // 2350
			  0 11101011 01010011011111001110110
	fp1 is = 1 11101010 10110011110110011101010,  -2.76253321865e+32
	fp2 is = 1 11101011 00101101011010011101011  -3.82086904847e+32


	fp1 is = 10100110011000110110001001001100, 	   -7.88896629161e-16
	fp2 is = 10101001100000011001010001010011,	   -5.7544809575e-14   ///847
	Error: expected = 0 01010010  11111111001101100011100, 
	     calculated = 0 01010010 11111111001101100011110

	Error: expected = 1 00001100 01000000111101011101010, /3171
	     calculated = 1 00001100 01000000111101011101100
	fp1 is = 0 00001001 01101010001000100001001, 
	fp2 is = 0 00001100 01101110001110100001100

	Error: expected = 0 11010001   10101011111011110101000, /3319
	     calculated = 0 11010011 01101010111110111101010
	fp1 is = 0 11010011 00111111011101111010011, 
	fp2 is = 0 11010010 10101000111101111010010
*/

/*
		temp_fraction = sol_frac[24:1];
		temp_exp = exp_in + 1'b1;

| (outallone == 1'b1)
 
Error: expected = 1 01010001 00001101010011101110001, 
     calculated = 1 01010000 11100101011000100011101

 	Error: expected = 1 11001000 10110101010000100000011, 
	     calculated = 1 11000110   00101010111101111110101
	fp1 is = 11100001001011001100111011000010,  -1.992336532e+20
	fp2 is = 01100100010101111110110111001000,  1.59327356825e+22

	Error: expected = 1 01010001 00001101010011101110001,  / 559
	     		  1 01010000  11100101011000100011100
				      0001101010011101110001111
	fp1 is = 1 01001110 01011000000111001001110,  -2.38775496161e-15
	fp2 is = 0 01010000 11000100100101101010000   1.25618509735e-14

	Error: expected = 1 01000111 00000001011011001101011, 
	     calculated = 1 01000110  11111101001001100101001   / 2143
	fp1 is = 1 01000100 01111010001111001000100,  -2.56302988134e-18
	fp2 is = 0 01000110 10100100010010101000110   1.13920157685e-17

	Error: expected = 1 10100111 01011001011000101111100, 
	     calculated = 1 10100110  01001101001110100000111  / 2437
	fp1 is = 1 10100101 10100101100111010100101,    -4.52705026048e+11
	fp2 is = 0 10100110 11011111111101110100110     1.03071914394e+12

	Error: expected = 1 10010010 00000101001101101010001, /  2450
	     calculated = 1 10010001  11110101100100101011101
	fp1 is = 1 10001110 10010111101100010001110,  -52184.5546875
	fp2 is = 0 10010001 11010111011101110010001   482780.53125

	Error: expected = 1 10100010 00000011010100010111010, /2626
	     calculated = 1 10100001  11111001010111010001011
	fp1 is = 1 10011110 11100000111111010011110,  -4034829824.0
	fp2 is = 0 10100001 11001010100000110100001   30770268160.0

	Error: expected = 1 11101100 00101101001110000110000, /2631
	     calculated = 1 11101011  10100101100011110100000	
	fp1 is = 1 11101010 00011001001100011101010,   -1.78228277794e+32
	fp2 is = 0 11101011 11001101110101111101011    5.85455694501e+32

	Error: expected = 1 11000010 00011101101110010010000,  /3687
	     calculated = 1 11000001  11000100100011011011110
	fp1 is = 11100000010001010100011011000000,  -5.68610415203e+19
	fp2 is = 01100000101110110001010111000001   1.07847146123e+20

	Error: expected = 1 10000010 00000100001000000101010,  /3911
	     calculated = 1 10000001  11110111101111110101011
	fp1 is = 10111110000001001101101001111100, -0.129739701748
	fp2 is = 01000000111111111111100110000001  7.99920701981

	Error: expected = 1 01000001 01011011101110000101111,  /4184
	     calculated = 1 01000000  01001000100011110100000
	fp1 is = 10011111110000000110111000111111,  -8.14975497991e-20
	fp2 is = 00100000011110111000000101000000   2.13032922138e-19

	Error: expected = 1 01100001 00101001001010011000111, /4393 
	     calculated = 1 01100000  10101101101011001110000
	fp1 is = 10101111101011111001100001011111,  -3.19405807359e-10
	fp2 is = 00110000010100010101110101100000   7.61664509241e-10

	Error: expected = 1 11011110 00001100100010110100101, /4464
	     calculated = 1 11011101  11100110111010010110101
	fp1 is = 1 11011100 00111000101001011011100, 
	fp2 is = 0 11011101 01111100110000111011101

	Error: expected = 1 11010011 01110100110100000011101, 
	     calculated = 1 11010010  00010110010111111000101

	Error: expected = 1 01100000 00111111100010101101101, 
	     calculated = 1 01100000 00111111100010101101100

	 Error: expected = 1 00101111 10101011111000001000110, 
	      calculated = 1 00101111 10101011111000001000101
*/


/*
	Error: expected = 1 11001000 10110101010000100000011, 
	     calculated = 1 11000110 00101010111101111110101,	
	fp1 is = 11100001001011001100111011000010,  -1.992336532e+20
	fp2 is = 01100100010101111110110111001000   1.59327356825e+22

	Error: expected = 1 11001000 10110101010000100000011, 
	     calculated = 1 11001000 01001010101111011111101

	Error: expected = 1 00011100 10000010100010100101011, 
	     calculated = 1 00011010 11110101110101101010011,
	fp1 is = 10000100011101111110010000001000,  -2.91394172802e-36
	fp2 is = 00001110010000010100010100011100   2.38223616268e-30
	
	Error: expected = 1 00011100 10000010100010100101011, 
	     calculated = 1 00011100 01111101011101011010100

	Error: expected = 1 01010001 00001101010011101110001, 
	     calculated = 1 01010000  00011010100111011100011,
	fp1 is = 10100111001011000000111001001110,  -2.38775496161e-15
	fp2 is = 00101000011000100100101101010000   1.25618509735e-14
*/

/*
Error: expected = 1 01010001 00001101010011101110001, -1.49496046645e-14
     calculated = 1 01010000  11100101011000100011101,  -1.34721039188e-14
wrong case =         559,
fp1 is = 1 01001110 01011000000111001001110,  -2.38775496161e-15
fp2 is = 0 01010000 11000100100101101010000, 1.25618509735e-14
 
Error: expected = 1 01000111 00000001011011001101011, -1.39550448227e-17
     calculated = 1 01000110  11111101001001100101001,  -1.38005299658e-17
wrong case =        2143,, 
fp1 is = 1 01000100 01111010001111001000100,  -2.56302988134e-18
fp2 is = 0 01000110 10100100010010101000110,  1.13920157685e-17

Error: expected = 1 10100111 01011001011000101111100, -1.48342413722e+12
     calculated = 1 10100110  01001101001110100001000, -7.15599118336e+11
wrong case =        2437,  
fp1 is = 1 10100101 10100101100111010100101, -4.52705026048e+11
fp2 is = 0 10100110 11011111111101110100110, 1.03071914394e+12

Error: expected = 1 10010010 00000101001101101010001, -534965.0625
     calculated = 1 10010001  11110101100100101011101,  -513610.90625
wrong case =        2450,
fp1 is = 1 10001110 10010111101100010001110, -52184.5546875
fp2 is = 0 10010001  11010111011101110010001, 482780.53125

Error: expected = 1 10100010 00000011010100010111010, -34805096448.0
     calculated = 1 10100001  11111001010111010001011, -33914378240.0
wrong case =        2626, 
fp1 is = 1 10011110 11100000111111010011110, -4034829824.0
fp2 is = 0 10100001 11001010100000110100001,  30770268160.0

Error: expected = 1 11101100 00101101001110000110000, -7.63683972295e+32
     calculated = 1 11101011  10100101100011110100000, -5.34390242339e+32
wrong case =        2631, , 
fp1 is = 1 11101010 00011001001100011101010,  -1.78228277794e+32
fp2 is = 0 11101011 11001101110101111101011,  5.85455694501e+32

Error: expected = 1 11000010 00011101101110010010000, -1.64708178847e+20
     calculated = 1 11000001  11000100100011011011111, -1.30439717536e+20
wrong case =        3687,  
fp1 is = 1 11000000 10001010100011011000000, -5.68610415203e+19
fp2 is = 0 11000001 01110110001010111000001, 1.07847146123e+20

Error: expected = 1 10000010 00000100001000000101010, -8.12894630432
     calculated = 1 10000001  11110111101111110101011, -7.87105321884
wrong case =        3911,  
fp1 is = 1 01111100 00001001101101001111100, -0.129739701748
fp2 is = 0 10000001 11111111111100110000001, 7.99920701981

Error: expected = 1 01000001 01011011101110000101111, -2.9453045255e-19
     calculated = 1 01000000  01001000100011110100000,  -1.39150390595e-19
wrong case =        4184, 
fp1 is = 1 00111111 10000000110111000111111,  -8.14975497991e-20
fp2 is = 0 01000000 11110111000000101000000,  2.13032922138e-19

Error: expected = 1 01100001 00101001001010011000111,  -1.08107023333e-09
     calculated = 1 01100000  10101101101011001110001,  -7.81574860387e-10
wrong case =        4393, 
fp1 is = 1 01011111 01011111001100001011111, -3.19405807359e-10
fp2 is = 0 01100000 10100010101110101100000, 7.61664509241e-10

Error: expected = 1 11011110 00001100100010110100101,  -4.15551863881e+28
     calculated = 1 11011101  11100110111010010110101,      -3.7672973765e+28
wrong case =        4464,  
fp1 is = 1 11011100 00111000101001011011100, -1.20949580925e+28
fp2 is = 0 11011101 01111100110000111011101,  2.94602306568e+28

Error: expected = 1 00100100 01000010000010000011010, -5.08076978623e-28
     calculated = 1 00100011  01111011111011111001011,  -2.99716564249e-28
wrong case =        4523,, 
fp1 is = 1 00100010 01111111000101000100010,  -1.51098087489e-28
fp2 is = 0 00100011 11000100100001100100011,  3.56978891134e-28

Error: expected = 1 11111100 00011100001000000111100,  -4.72086672739e+37
     calculated = 1 11111011  11000111101111110001000,  -3.78619244563e+37
wrong case =        4720,
fp1 is = 1 11111010 10010000000010011111010,  -1.66169649342e+37
fp2 is = 0 11111011 01110000001110111111011,  3.05917023398e+37

Error: expected = 1 10010100 01000111100111101101110,  -2683867.5
     calculated = 1 10010011  01110000110000100100011,  -1510436.375
wrong case =        4941,  
fp1 is = 1 10010010 00110001111111010010010, -626665.125
fp2 is = 0 10010011 11110110001111110010011, 2057202.375

Error: expected = 1 01111010 00000111001010001011010,  -0.03212390095
     calculated = 1 01111001  111110001101011101001011,   -0.0303760971874
wrong case =        5210,  
fp1 is = 1 01111000 11111111100111001111000,  -0.0156131908298
fp2 is = 0 01111001 00001110100000101111001,  0.0165107119828

Error: expected = 1 01100110 00001100010011100111110,  -3.12349968112e-08
     calculated = 1 01100101  11100111011000110000010,  -2.83696444114e-08
wrong case =        5262, 
fp1 is = 1 01100011 10110101010110001100011,  -6.36423314049e-09
fp2 is = 0 01100101 10101011010001101100101,  2.48707667794e-08
 
Error: expected = 1 00100111 00010000010100010011100, -3.43712705306e-27
     calculated = 1 00100110  11011111010111011000111, -3.02522128992e-27
wrong case =        6621,  
fp1 is = 1 00100101 00101111111100000100101,  -9.59061208493e-28
fp2 is = 0 00100110 10001000101010100100110,  2.47806594087e-27

Error: expected = 1 00111100 00110101110011100101100,  -8.20049734061e-21
     calculated = 1 00111011  10010100011000110101000, -5.35202981545e-21
wrong case =        7260,  
fp1 is = 1 00111010 10010000111111000111010,  -2.6535037205e-21
fp2 is = 0 00111011 10100011000111100111011,  5.54699362011e-21

Error: expected = 1 10001000 01101100000110101100101,  -728.209289551
     calculated = 1 10000111 00100111110010100110101,  -295.790679932
wrong case =        8721,  
fp1 is = 1 10000110 11110110111011010000110,  -251.462982178
fp2 is = 0 10000111 11011100101111110000111,  476.746307373

Error: expected = 1 10100101 00010111000101111111010,  -2.99674435584e+11
     calculated = 1 10100100 11010001110100000001011,  -2.5008136192e+11
wrong case =        9087,  
fp1 is = 1 10100011 11100011110110010100011, -1.2988215296e+11
fp2 is = 0 10100100 00111100010000110100100, 1.697923072e+11

Error: expected = 1 00001100 00001011001011100001000, -2.51254800237e-35
     calculated = 1 00001011  11101001101000111110000,  -2.30227685859e-35
wrong case =        9225,  
fp1 is = 1 00001010 10010101000001000001010, -9.52187875829e-36
fp2 is = 0 00001011 01001011110110100001011,  1.56036012654e-35

Error: expected = 1 11010011 01110100110100000011101, -2.81689829398e+25
     calculated = 1 11010010  00010110010111111000101,  -1.0516642135e+25
wrong case =        9954,
fp1 is = 1 11010001 11111000000110011010001,  -9.52218219719e+24
fp2 is = 0 11010010 11101101100100111010010,  1.8646801319e+25




Error: expected = 10110110001000000000000000000000, calculated = 10110110000000000010100000000000, wrong case =        6655,  fp1 is = 00111100000110101100000101111000, fp2 is = 00111100000110101100101101111000, 
*/


/*
Error: expected = 1 00000100 11111101100000010000100,-1.87162220941e-37
     calculated = 1 00000000 00000000000000000000000, -0.0
wrong case =      146985,  
fp1 is = 1 00000000 10011010101100000000000, -7.10290165597e-39
fp2 is = 0 00000100 11100011110101100000100, 1.77733298359e-37

Error: expected = 1 00001011 11111111111100100001101, -2.4071571565e-35
     calculated = 1 00000000 00000000000000000000000,  -0.0
wrong case =      161537,  
fp1 is = 1 00001001 01100101011000000001001,  -4.20092616484e-36
fp2 is = 0 00001011 10100110100110100001011, 1.98706457589e-35

Error: expected = 10000011011111100101110100010110, -7.47507486929e-37
     calculated = 10000000000000000000000000000000, -0.0
wrong case =      198397,
fp1 is = 1 00000000 11001100000010000000000,  -9.36865553774e-39
fp2 is = 0 00000110 11110101100010100000110,  7.36945687406e-37


*/

	 if(floating_point1[30:23] == 8'b11111111) 
	   floating_point1[30:23] = 8'b11111110;
	 if(floating_point2[30:23] == 8'b11111111) 
	   floating_point2[30:23] = 8'b11111110;

	 //convert from floating point to 2 real values
	 fp_convert(.val(floating_point1), .fp(fp1_real));
	 fp_convert(.val(floating_point2), .fp(fp2_real));

	 //performing real number arithemetic
	 //
	 if(funct7 == 7'b0100000) begin
	    result_real = fp1_real + fp2_real; //addition
	 end else if (funct7 == 7'b0000010) begin
	    result_real = fp1_real * fp2_real; //multiplication
         end else if (funct7 == 7'b0100100) begin
	    result_real = fp1_real - fp2_real; //subtraction
	 end
	 
	 else result_real = 'x;
	 
	 real_to_fp(.r(result_real), .fp(result_binary)); //convert the real number back to floating point
	 @(negedge clk);
	 @(negedge clk);
	 fp_convert(.val(floating_point_out), .fp(fp_out_real));
	 #1;
	 assert((floating_point_out == result_binary) || (floating_point_out == result_binary + 1)) 
	   else begin
	      j = j + 1;
	      $error("expected = %b, calculated = %b, wrong case = %d, number = %d, fp1 is = %b, fp2 is = %b, result_real is %d", result_binary, floating_point_out, i, j, floating_point1, floating_point2, result_real);
	//$error("expected = %b, calculated = %b, wrong case = %d, number = %d", result_binary, floating_point_out, i, j);
	      //$display(fp1_real);//
	      //$display(fp2_real);//
	      //$display(result_real); //expected
	      //$display(fp_out_real); //computed
	   end
	 //if((flags[1] == 0) & (flags[2] == 0)) begin
	   // assert(flags[0] == 0) else $error("asdklfj;as");
	 //end
	 @(negedge clk);
	 floating_point1 = 'x;
	 floating_point2 = 'x;
	 frm             = 'x;
	 funct7          = 'x;
	 result_real     = 'x;
	 fp1_real        = 'x;
	 fp2_real        = 'x;
	 fp_exp          = 'x;
	 fp_frac         = 'x;
	 @(negedge clk);
	 
      end
   endtask // random_check
   
   task real_to_fp;
      input shortreal r;
      output reg [31:0] fp;
      begin
	 
	 int fp_index;
	 shortreal MAX;
	 shortreal MIN;
	 
	 fp_convert(32'b01111111011111111111111111111111, MAX);
	 fp_convert(32'b00000000000000000000000000000000, MIN);
	 
	 
	 fp = 32'b01000000000000000000000000000000;

	 if(r < 0) begin // set sign bit
	    fp[31] = 1'b1;
	    r = -r;
	 end
	 
	 if(r < MIN) // ovf 
	    fp[30:0] = 31'b0000000000000000000000000000000;
	 
         else if(r > MAX) // unf
	    fp[30:0] = 31'b1111111100000000000000000000000;
	 
	 else begin // everything else
	    if(r >= 2) begin 
	       while(r >= 2) begin
	          r /= 2;
		  fp[30:23] += 1;
	       end
	    end
	    else if(r < 1) begin
	       while(r < 1) begin
		  r *= 2;
		  fp[30:23] -= 1;
	       end
	    end
	    
	    r -= 1;
	    fp_index = 22;
	    for(shortreal i = 0.50; i != 2**-24; i /= 2) begin
	       if(r >= i) begin
		  r -= i;
		  fp[fp_index] = 1'b1;
	       end
	       fp_index -= 1;
	    end
	 end // else: !if((r>(1.70141*(10**38))))
      end
   endtask // real_to_fp
         
   task fp_convert;
      input [31:0] val;
      output shortreal  fp;
      begin
         
	 fp_exp  = shortreal'(val[30:23]);
	 fp_frac = shortreal'(val[22:0]);

	 fp_exp = fp_exp - 128;
	 
	 for(int k = 0; k < 23; k = k + 1) begin
	    fp_frac /= 2;
	 end
     	 fp_frac = fp_frac + 1;	 

	 if(val[31]) 
	   fp = -fp_frac * (2 ** fp_exp);
	 else
	   fp = fp_frac * (2 ** fp_exp);
      end
   endtask // fp_convert
   
initial begin
   nrst = 1;
   @(negedge clk);
   nrst = 0;
   @(negedge clk);
   nrst = 1;
   i = 0;

   /*while((i <= 62))begin
      random_check();
      i = i + 1;
      //break;
      end //*/
   while (1) begin
	i = i + 1;
	random_check();
  end //*/
end
   
endmodule // tb_FPU_top_level
