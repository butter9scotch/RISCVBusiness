`ifndef RV32V_LOADSTORE_UNIT_IF_VH
`define RV32V_LOADSTORE_UNIT_IF_VH

interface rv32v_loadstore_unit_if();



endinterface

`endif //RV32V_LOADSTORE_UNIT_IF_VH