module rv32v_top_level();


  
endmodule