module add_unsigned_GENERIC_REAL(A, B, Z);
// synthesis_equation add_unsigned
  input [26:0] A, B;
  output [26:0] Z;
  wire [26:0] A, B;
  wire [26:0] Z;
  wire n_83, n_86, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_96, n_97, n_98, n_99, n_100, n_102, n_103, n_104;
  wire n_105, n_106, n_108, n_109, n_110, n_111, n_112, n_114;
  wire n_115, n_116, n_117, n_118, n_120, n_121, n_122, n_123;
  wire n_124, n_126, n_127, n_128, n_129, n_130, n_132, n_133;
  wire n_134, n_135, n_136, n_138, n_139, n_140, n_141, n_142;
  wire n_144, n_145, n_146, n_147, n_148, n_150, n_151, n_152;
  wire n_153, n_154, n_156, n_157, n_158, n_159, n_160, n_162;
  wire n_163, n_165, n_166, n_167, n_168, n_169, n_170, n_172;
  wire n_174, n_176, n_177, n_179, n_180, n_182, n_184, n_186;
  wire n_187, n_189, n_190, n_192, n_194, n_196, n_197, n_199;
  wire n_200, n_202, n_204, n_206, n_207, n_209, n_210, n_212;
  wire n_214, n_216, n_217, n_219, n_220, n_221, n_224, n_226;
  wire n_228, n_229, n_230, n_232, n_233, n_234, n_236, n_237;
  wire n_238, n_239, n_241, n_243, n_245, n_246, n_247, n_249;
  wire n_250, n_251, n_253, n_254, n_256, n_258, n_260, n_261;
  wire n_262, n_264, n_265, n_266, n_268, n_270, n_271, n_272;
  wire n_274, n_275, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_293, n_296, n_303, n_305, n_306, n_307, n_309;
  wire n_310, n_312, n_313, n_314, n_315, n_316, n_317, n_318;
  wire n_319, n_320, n_321, n_322, n_323, n_325, n_326, n_327;
  wire n_329, n_330, n_335, n_336, n_338, n_339, n_340, n_342;
  wire n_343, n_344, n_345, n_347, n_348, n_349, n_351, n_352;
  wire n_353, n_354, n_356, n_357, n_359, n_360, n_362, n_363;
  wire n_364, n_365, n_367, n_368, n_369, n_371, n_372, n_373;
  wire n_374, n_376, n_377, n_379, n_380, n_382, n_383, n_384;
  wire n_385, n_387, n_388, n_389, n_390, n_392, n_393, n_394;
  wire n_395;
  xor g1 (Z[0], A[0], B[0]);
  nand g2 (n_83, A[0], B[0]);
  nor g6 (n_86, A[1], B[1]);
  nand g7 (n_89, A[1], B[1]);
  nor g8 (n_96, A[2], B[2]);
  nand g9 (n_91, A[2], B[2]);
  nor g10 (n_92, A[3], B[3]);
  nand g11 (n_93, A[3], B[3]);
  nor g12 (n_102, A[4], B[4]);
  nand g13 (n_97, A[4], B[4]);
  nor g14 (n_98, A[5], B[5]);
  nand g15 (n_99, A[5], B[5]);
  nor g16 (n_108, A[6], B[6]);
  nand g17 (n_103, A[6], B[6]);
  nor g18 (n_104, A[7], B[7]);
  nand g19 (n_105, A[7], B[7]);
  nor g20 (n_114, A[8], B[8]);
  nand g21 (n_109, A[8], B[8]);
  nor g22 (n_110, A[9], B[9]);
  nand g23 (n_111, A[9], B[9]);
  nor g24 (n_120, A[10], B[10]);
  nand g25 (n_115, A[10], B[10]);
  nor g26 (n_116, A[11], B[11]);
  nand g27 (n_117, A[11], B[11]);
  nor g28 (n_126, A[12], B[12]);
  nand g29 (n_121, A[12], B[12]);
  nor g30 (n_122, A[13], B[13]);
  nand g31 (n_123, A[13], B[13]);
  nor g32 (n_132, A[14], B[14]);
  nand g33 (n_127, A[14], B[14]);
  nor g34 (n_128, A[15], B[15]);
  nand g35 (n_129, A[15], B[15]);
  nor g36 (n_138, A[16], B[16]);
  nand g37 (n_133, A[16], B[16]);
  nor g38 (n_134, A[17], B[17]);
  nand g39 (n_135, A[17], B[17]);
  nor g40 (n_144, A[18], B[18]);
  nand g41 (n_139, A[18], B[18]);
  nor g42 (n_140, A[19], B[19]);
  nand g43 (n_141, A[19], B[19]);
  nor g44 (n_150, A[20], B[20]);
  nand g45 (n_145, A[20], B[20]);
  nor g46 (n_146, A[21], B[21]);
  nand g47 (n_147, A[21], B[21]);
  nor g48 (n_156, A[22], B[22]);
  nand g49 (n_151, A[22], B[22]);
  nor g50 (n_152, A[23], B[23]);
  nand g51 (n_153, A[23], B[23]);
  nor g52 (n_162, A[24], B[24]);
  nand g53 (n_157, A[24], B[24]);
  nor g54 (n_158, A[25], B[25]);
  nand g55 (n_159, A[25], B[25]);
  nor g56 (n_219, A[26], B[26]);
  nand g57 (n_221, A[26], B[26]);
  nand g60 (n_163, n_89, n_90);
  nor g61 (n_94, n_91, n_92);
  nor g64 (n_166, n_96, n_92);
  nor g65 (n_100, n_97, n_98);
  nor g68 (n_172, n_102, n_98);
  nor g69 (n_106, n_103, n_104);
  nor g72 (n_174, n_108, n_104);
  nor g73 (n_112, n_109, n_110);
  nor g76 (n_182, n_114, n_110);
  nor g77 (n_118, n_115, n_116);
  nor g80 (n_184, n_120, n_116);
  nor g81 (n_124, n_121, n_122);
  nor g84 (n_192, n_126, n_122);
  nor g85 (n_130, n_127, n_128);
  nor g88 (n_194, n_132, n_128);
  nor g89 (n_136, n_133, n_134);
  nor g92 (n_202, n_138, n_134);
  nor g93 (n_142, n_139, n_140);
  nor g96 (n_204, n_144, n_140);
  nor g97 (n_148, n_145, n_146);
  nor g100 (n_212, n_150, n_146);
  nor g101 (n_154, n_151, n_152);
  nor g104 (n_214, n_156, n_152);
  nor g105 (n_160, n_157, n_158);
  nor g108 (n_224, n_162, n_158);
  nand g111 (n_338, n_91, n_165);
  nand g112 (n_168, n_166, n_163);
  nand g113 (n_226, n_167, n_168);
  nor g114 (n_170, n_108, n_169);
  nand g123 (n_234, n_172, n_174);
  nor g124 (n_180, n_120, n_179);
  nand g133 (n_241, n_182, n_184);
  nor g134 (n_190, n_132, n_189);
  nand g143 (n_249, n_192, n_194);
  nor g144 (n_200, n_144, n_199);
  nand g153 (n_256, n_202, n_204);
  nor g154 (n_210, n_156, n_209);
  nand g163 (n_264, n_212, n_214);
  nand g171 (n_342, n_97, n_228);
  nand g172 (n_229, n_172, n_226);
  nand g173 (n_344, n_169, n_229);
  nand g176 (n_347, n_232, n_233);
  nand g179 (n_268, n_236, n_237);
  nor g180 (n_239, n_126, n_238);
  nor g183 (n_278, n_126, n_241);
  nor g189 (n_247, n_245, n_238);
  nor g192 (n_284, n_241, n_245);
  nor g193 (n_251, n_249, n_238);
  nor g196 (n_287, n_241, n_249);
  nor g197 (n_254, n_150, n_253);
  nor g200 (n_313, n_150, n_256);
  nor g206 (n_262, n_260, n_253);
  nor g209 (n_319, n_256, n_260);
  nor g210 (n_266, n_264, n_253);
  nor g213 (n_293, n_256, n_264);
  nand g216 (n_351, n_109, n_270);
  nand g217 (n_271, n_182, n_268);
  nand g218 (n_353, n_179, n_271);
  nand g221 (n_356, n_274, n_275);
  nand g224 (n_359, n_238, n_277);
  nand g225 (n_280, n_278, n_268);
  nand g226 (n_362, n_279, n_280);
  nand g227 (n_283, n_281, n_268);
  nand g228 (n_364, n_282, n_283);
  nand g229 (n_286, n_284, n_268);
  nand g230 (n_367, n_285, n_286);
  nand g231 (n_289, n_287, n_268);
  nand g232 (n_303, n_288, n_289);
  nor g233 (n_291, n_162, n_290);
  nand g242 (n_327, n_224, n_293);
  nand g250 (n_371, n_133, n_305);
  nand g251 (n_306, n_202, n_303);
  nand g252 (n_373, n_199, n_306);
  nand g255 (n_376, n_309, n_310);
  nand g258 (n_379, n_253, n_312);
  nand g259 (n_315, n_313, n_303);
  nand g260 (n_382, n_314, n_315);
  nand g261 (n_318, n_316, n_303);
  nand g262 (n_384, n_317, n_318);
  nand g263 (n_321, n_319, n_303);
  nand g264 (n_387, n_320, n_321);
  nand g265 (n_322, n_293, n_303);
  nand g266 (n_389, n_290, n_322);
  nand g269 (n_392, n_325, n_326);
  nand g272 (n_394, n_329, n_330);
  xnor g279 (Z[2], n_163, n_336);
  xnor g282 (Z[3], n_338, n_339);
  xnor g284 (Z[4], n_226, n_340);
  xnor g287 (Z[5], n_342, n_343);
  xnor g289 (Z[6], n_344, n_345);
  xnor g292 (Z[7], n_347, n_348);
  xnor g294 (Z[8], n_268, n_349);
  xnor g297 (Z[9], n_351, n_352);
  xnor g299 (Z[10], n_353, n_354);
  xnor g302 (Z[11], n_356, n_357);
  xnor g305 (Z[12], n_359, n_360);
  xnor g308 (Z[13], n_362, n_363);
  xnor g310 (Z[14], n_364, n_365);
  xnor g313 (Z[15], n_367, n_368);
  xnor g315 (Z[16], n_303, n_369);
  xnor g318 (Z[17], n_371, n_372);
  xnor g320 (Z[18], n_373, n_374);
  xnor g323 (Z[19], n_376, n_377);
  xnor g326 (Z[20], n_379, n_380);
  xnor g329 (Z[21], n_382, n_383);
  xnor g331 (Z[22], n_384, n_385);
  xnor g334 (Z[23], n_387, n_388);
  xnor g336 (Z[24], n_389, n_390);
  xnor g339 (Z[25], n_392, n_393);
  xnor g341 (Z[26], n_394, n_395);
  or g344 (n_90, n_83, n_86);
  and g345 (n_167, wc, n_93);
  not gc (wc, n_94);
  and g346 (n_169, wc0, n_99);
  not gc0 (wc0, n_100);
  and g347 (n_176, wc1, n_105);
  not gc1 (wc1, n_106);
  and g348 (n_179, wc2, n_111);
  not gc2 (wc2, n_112);
  and g349 (n_186, wc3, n_117);
  not gc3 (wc3, n_118);
  and g350 (n_189, wc4, n_123);
  not gc4 (wc4, n_124);
  and g351 (n_196, wc5, n_129);
  not gc5 (wc5, n_130);
  and g352 (n_199, wc6, n_135);
  not gc6 (wc6, n_136);
  and g353 (n_206, wc7, n_141);
  not gc7 (wc7, n_142);
  and g354 (n_209, wc8, n_147);
  not gc8 (wc8, n_148);
  and g355 (n_216, wc9, n_153);
  not gc9 (wc9, n_154);
  and g356 (n_220, wc10, n_159);
  not gc10 (wc10, n_160);
  or g357 (n_230, wc11, n_108);
  not gc11 (wc11, n_172);
  or g358 (n_272, wc12, n_120);
  not gc12 (wc12, n_182);
  or g359 (n_245, wc13, n_132);
  not gc13 (wc13, n_192);
  or g360 (n_307, wc14, n_144);
  not gc14 (wc14, n_202);
  or g361 (n_260, wc15, n_156);
  not gc15 (wc15, n_212);
  or g362 (n_335, wc16, n_86);
  not gc16 (wc16, n_89);
  or g363 (n_336, wc17, n_96);
  not gc17 (wc17, n_91);
  or g364 (n_339, wc18, n_92);
  not gc18 (wc18, n_93);
  or g365 (n_340, wc19, n_102);
  not gc19 (wc19, n_97);
  or g366 (n_343, wc20, n_98);
  not gc20 (wc20, n_99);
  or g367 (n_345, wc21, n_108);
  not gc21 (wc21, n_103);
  or g368 (n_348, wc22, n_104);
  not gc22 (wc22, n_105);
  or g369 (n_349, wc23, n_114);
  not gc23 (wc23, n_109);
  or g370 (n_352, wc24, n_110);
  not gc24 (wc24, n_111);
  or g371 (n_354, wc25, n_120);
  not gc25 (wc25, n_115);
  or g372 (n_357, wc26, n_116);
  not gc26 (wc26, n_117);
  or g373 (n_360, wc27, n_126);
  not gc27 (wc27, n_121);
  or g374 (n_363, wc28, n_122);
  not gc28 (wc28, n_123);
  or g375 (n_365, wc29, n_132);
  not gc29 (wc29, n_127);
  or g376 (n_368, wc30, n_128);
  not gc30 (wc30, n_129);
  or g377 (n_369, wc31, n_138);
  not gc31 (wc31, n_133);
  or g378 (n_372, wc32, n_134);
  not gc32 (wc32, n_135);
  or g379 (n_374, wc33, n_144);
  not gc33 (wc33, n_139);
  or g380 (n_377, wc34, n_140);
  not gc34 (wc34, n_141);
  or g381 (n_380, wc35, n_150);
  not gc35 (wc35, n_145);
  or g382 (n_383, wc36, n_146);
  not gc36 (wc36, n_147);
  or g383 (n_385, wc37, n_156);
  not gc37 (wc37, n_151);
  or g384 (n_388, wc38, n_152);
  not gc38 (wc38, n_153);
  or g385 (n_390, wc39, n_162);
  not gc39 (wc39, n_157);
  or g386 (n_393, wc40, n_158);
  not gc40 (wc40, n_159);
  or g387 (n_395, wc41, n_219);
  not gc41 (wc41, n_221);
  and g388 (n_177, wc42, n_174);
  not gc42 (wc42, n_169);
  and g389 (n_187, wc43, n_184);
  not gc43 (wc43, n_179);
  and g390 (n_197, wc44, n_194);
  not gc44 (wc44, n_189);
  and g391 (n_207, wc45, n_204);
  not gc45 (wc45, n_199);
  and g392 (n_217, wc46, n_214);
  not gc46 (wc46, n_209);
  and g393 (n_281, wc47, n_192);
  not gc47 (wc47, n_241);
  and g394 (n_316, wc48, n_212);
  not gc48 (wc48, n_256);
  xor g395 (Z[1], n_83, n_335);
  or g396 (n_165, wc49, n_96);
  not gc49 (wc49, n_163);
  and g397 (n_232, wc50, n_103);
  not gc50 (wc50, n_170);
  and g398 (n_236, wc51, n_176);
  not gc51 (wc51, n_177);
  and g399 (n_274, wc52, n_115);
  not gc52 (wc52, n_180);
  and g400 (n_238, wc53, n_186);
  not gc53 (wc53, n_187);
  and g401 (n_246, wc54, n_127);
  not gc54 (wc54, n_190);
  and g402 (n_250, wc55, n_196);
  not gc55 (wc55, n_197);
  and g403 (n_309, wc56, n_139);
  not gc56 (wc56, n_200);
  and g404 (n_253, wc57, n_206);
  not gc57 (wc57, n_207);
  and g405 (n_261, wc58, n_151);
  not gc58 (wc58, n_210);
  and g406 (n_265, wc59, n_216);
  not gc59 (wc59, n_217);
  or g407 (n_323, wc60, n_162);
  not gc60 (wc60, n_293);
  and g408 (n_243, wc61, n_192);
  not gc61 (wc61, n_238);
  and g409 (n_258, wc62, n_212);
  not gc62 (wc62, n_253);
  or g410 (n_228, wc63, n_102);
  not gc63 (wc63, n_226);
  or g411 (n_233, n_230, wc64);
  not gc64 (wc64, n_226);
  or g412 (n_237, n_234, wc65);
  not gc65 (wc65, n_226);
  and g413 (n_279, wc66, n_121);
  not gc66 (wc66, n_239);
  and g414 (n_282, wc67, n_189);
  not gc67 (wc67, n_243);
  and g415 (n_285, n_246, wc68);
  not gc68 (wc68, n_247);
  and g416 (n_288, n_250, wc69);
  not gc69 (wc69, n_251);
  and g417 (n_314, wc70, n_145);
  not gc70 (wc70, n_254);
  and g418 (n_317, wc71, n_209);
  not gc71 (wc71, n_258);
  and g419 (n_320, n_261, wc72);
  not gc72 (wc72, n_262);
  and g420 (n_290, n_265, wc73);
  not gc73 (wc73, n_266);
  and g421 (n_296, wc74, n_224);
  not gc74 (wc74, n_290);
  or g422 (n_270, wc75, n_114);
  not gc75 (wc75, n_268);
  or g423 (n_275, n_272, wc76);
  not gc76 (wc76, n_268);
  or g424 (n_277, wc77, n_241);
  not gc77 (wc77, n_268);
  and g425 (n_325, wc78, n_157);
  not gc78 (wc78, n_291);
  and g426 (n_329, wc79, n_220);
  not gc79 (wc79, n_296);
  or g427 (n_305, wc80, n_138);
  not gc80 (wc80, n_303);
  or g428 (n_310, n_307, wc81);
  not gc81 (wc81, n_303);
  or g429 (n_312, wc82, n_256);
  not gc82 (wc82, n_303);
  or g430 (n_326, n_323, wc83);
  not gc83 (wc83, n_303);
  or g431 (n_330, n_327, wc84);
  not gc84 (wc84, n_303);
endmodule

module add_unsigned_GENERIC(A, B, Z);
  input [26:0] A, B;
  output [26:0] Z;
  wire [26:0] A, B;
  wire [26:0] Z;
  add_unsigned_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

