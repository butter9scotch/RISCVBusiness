module add_unsigned_GENERIC_REAL(A, B, Z);
// synthesis_equation add_unsigned
  input [26:0] A, B;
  output [26:0] Z;
  wire [26:0] A, B;
  wire [26:0] Z;
  wire n_83, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190;
  wire n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198;
  wire n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_207, n_208, n_209, n_210, n_211, n_212, n_216;
  nand g1 (n_83, A[0], B[0]);
  xor g5 (Z[0], A[0], B[0]);
  nand g7 (n_88, A[1], B[1]);
  nand g10 (n_92, n_88, n_89, n_90);
  xor g11 (n_91, A[1], B[1]);
  nand g13 (n_93, A[2], B[2]);
  nand g14 (n_94, A[2], n_92);
  nand g15 (n_95, B[2], n_92);
  nand g16 (n_97, n_93, n_94, n_95);
  xor g17 (n_96, A[2], B[2]);
  xor g18 (Z[2], n_92, n_96);
  nand g19 (n_98, A[3], B[3]);
  nand g20 (n_99, A[3], n_97);
  nand g21 (n_100, B[3], n_97);
  nand g22 (n_102, n_98, n_99, n_100);
  xor g23 (n_101, A[3], B[3]);
  xor g24 (Z[3], n_97, n_101);
  nand g25 (n_103, A[4], B[4]);
  nand g26 (n_104, A[4], n_102);
  nand g27 (n_105, B[4], n_102);
  nand g28 (n_107, n_103, n_104, n_105);
  xor g29 (n_106, A[4], B[4]);
  xor g30 (Z[4], n_102, n_106);
  nand g31 (n_108, A[5], B[5]);
  nand g32 (n_109, A[5], n_107);
  nand g33 (n_110, B[5], n_107);
  nand g34 (n_112, n_108, n_109, n_110);
  xor g35 (n_111, A[5], B[5]);
  xor g36 (Z[5], n_107, n_111);
  nand g37 (n_113, A[6], B[6]);
  nand g38 (n_114, A[6], n_112);
  nand g39 (n_115, B[6], n_112);
  nand g40 (n_117, n_113, n_114, n_115);
  xor g41 (n_116, A[6], B[6]);
  xor g42 (Z[6], n_112, n_116);
  nand g43 (n_118, A[7], B[7]);
  nand g44 (n_119, A[7], n_117);
  nand g45 (n_120, B[7], n_117);
  nand g46 (n_122, n_118, n_119, n_120);
  xor g47 (n_121, A[7], B[7]);
  xor g48 (Z[7], n_117, n_121);
  nand g49 (n_123, A[8], B[8]);
  nand g50 (n_124, A[8], n_122);
  nand g51 (n_125, B[8], n_122);
  nand g52 (n_127, n_123, n_124, n_125);
  xor g53 (n_126, A[8], B[8]);
  xor g54 (Z[8], n_122, n_126);
  nand g55 (n_128, A[9], B[9]);
  nand g56 (n_129, A[9], n_127);
  nand g57 (n_130, B[9], n_127);
  nand g58 (n_132, n_128, n_129, n_130);
  xor g59 (n_131, A[9], B[9]);
  xor g60 (Z[9], n_127, n_131);
  nand g61 (n_133, A[10], B[10]);
  nand g62 (n_134, A[10], n_132);
  nand g63 (n_135, B[10], n_132);
  nand g64 (n_137, n_133, n_134, n_135);
  xor g65 (n_136, A[10], B[10]);
  xor g66 (Z[10], n_132, n_136);
  nand g67 (n_138, A[11], B[11]);
  nand g68 (n_139, A[11], n_137);
  nand g69 (n_140, B[11], n_137);
  nand g70 (n_142, n_138, n_139, n_140);
  xor g71 (n_141, A[11], B[11]);
  xor g72 (Z[11], n_137, n_141);
  nand g73 (n_143, A[12], B[12]);
  nand g74 (n_144, A[12], n_142);
  nand g75 (n_145, B[12], n_142);
  nand g76 (n_147, n_143, n_144, n_145);
  xor g77 (n_146, A[12], B[12]);
  xor g78 (Z[12], n_142, n_146);
  nand g79 (n_148, A[13], B[13]);
  nand g80 (n_149, A[13], n_147);
  nand g81 (n_150, B[13], n_147);
  nand g82 (n_152, n_148, n_149, n_150);
  xor g83 (n_151, A[13], B[13]);
  xor g84 (Z[13], n_147, n_151);
  nand g85 (n_153, A[14], B[14]);
  nand g86 (n_154, A[14], n_152);
  nand g87 (n_155, B[14], n_152);
  nand g88 (n_157, n_153, n_154, n_155);
  xor g89 (n_156, A[14], B[14]);
  xor g90 (Z[14], n_152, n_156);
  nand g91 (n_158, A[15], B[15]);
  nand g92 (n_159, A[15], n_157);
  nand g93 (n_160, B[15], n_157);
  nand g94 (n_162, n_158, n_159, n_160);
  xor g95 (n_161, A[15], B[15]);
  xor g96 (Z[15], n_157, n_161);
  nand g97 (n_163, A[16], B[16]);
  nand g98 (n_164, A[16], n_162);
  nand g99 (n_165, B[16], n_162);
  nand g100 (n_167, n_163, n_164, n_165);
  xor g101 (n_166, A[16], B[16]);
  xor g102 (Z[16], n_162, n_166);
  nand g103 (n_168, A[17], B[17]);
  nand g104 (n_169, A[17], n_167);
  nand g105 (n_170, B[17], n_167);
  nand g106 (n_172, n_168, n_169, n_170);
  xor g107 (n_171, A[17], B[17]);
  xor g108 (Z[17], n_167, n_171);
  nand g109 (n_173, A[18], B[18]);
  nand g110 (n_174, A[18], n_172);
  nand g111 (n_175, B[18], n_172);
  nand g112 (n_177, n_173, n_174, n_175);
  xor g113 (n_176, A[18], B[18]);
  xor g114 (Z[18], n_172, n_176);
  nand g115 (n_178, A[19], B[19]);
  nand g116 (n_179, A[19], n_177);
  nand g117 (n_180, B[19], n_177);
  nand g118 (n_182, n_178, n_179, n_180);
  xor g119 (n_181, A[19], B[19]);
  xor g120 (Z[19], n_177, n_181);
  nand g121 (n_183, A[20], B[20]);
  nand g122 (n_184, A[20], n_182);
  nand g123 (n_185, B[20], n_182);
  nand g124 (n_187, n_183, n_184, n_185);
  xor g125 (n_186, A[20], B[20]);
  xor g126 (Z[20], n_182, n_186);
  nand g127 (n_188, A[21], B[21]);
  nand g128 (n_189, A[21], n_187);
  nand g129 (n_190, B[21], n_187);
  nand g130 (n_192, n_188, n_189, n_190);
  xor g131 (n_191, A[21], B[21]);
  xor g132 (Z[21], n_187, n_191);
  nand g133 (n_193, A[22], B[22]);
  nand g134 (n_194, A[22], n_192);
  nand g135 (n_195, B[22], n_192);
  nand g136 (n_197, n_193, n_194, n_195);
  xor g137 (n_196, A[22], B[22]);
  xor g138 (Z[22], n_192, n_196);
  nand g139 (n_198, A[23], B[23]);
  nand g140 (n_199, A[23], n_197);
  nand g141 (n_200, B[23], n_197);
  nand g142 (n_202, n_198, n_199, n_200);
  xor g143 (n_201, A[23], B[23]);
  xor g144 (Z[23], n_197, n_201);
  nand g145 (n_203, A[24], B[24]);
  nand g146 (n_204, A[24], n_202);
  nand g147 (n_205, B[24], n_202);
  nand g148 (n_207, n_203, n_204, n_205);
  xor g149 (n_206, A[24], B[24]);
  xor g150 (Z[24], n_202, n_206);
  nand g151 (n_208, A[25], B[25]);
  nand g152 (n_209, A[25], n_207);
  nand g153 (n_210, B[25], n_207);
  nand g154 (n_212, n_208, n_209, n_210);
  xor g155 (n_211, A[25], B[25]);
  xor g156 (Z[25], n_207, n_211);
  xor g161 (n_216, A[26], B[26]);
  xor g162 (Z[26], n_212, n_216);
  or g164 (n_89, wc, n_83);
  not gc (wc, A[1]);
  or g165 (n_90, wc0, n_83);
  not gc0 (wc0, B[1]);
  xnor g166 (Z[1], n_83, n_91);
endmodule

module add_unsigned_GENERIC(A, B, Z);
  input [26:0] A, B;
  output [26:0] Z;
  wire [26:0] A, B;
  wire [26:0] Z;
  add_unsigned_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_unsigned_161_GENERIC_REAL(A, B, Z);
// synthesis_equation add_unsigned
  input [26:0] A, B;
  output [26:0] Z;
  wire [26:0] A, B;
  wire [26:0] Z;
  wire n_83, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190;
  wire n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198;
  wire n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_207, n_208, n_209, n_210, n_211, n_212, n_216;
  nand g1 (n_83, A[0], B[0]);
  xor g5 (Z[0], A[0], B[0]);
  nand g7 (n_88, A[1], B[1]);
  nand g10 (n_92, n_88, n_89, n_90);
  xor g11 (n_91, A[1], B[1]);
  nand g13 (n_93, A[2], B[2]);
  nand g14 (n_94, A[2], n_92);
  nand g15 (n_95, B[2], n_92);
  nand g16 (n_97, n_93, n_94, n_95);
  xor g17 (n_96, A[2], B[2]);
  xor g18 (Z[2], n_92, n_96);
  nand g19 (n_98, A[3], B[3]);
  nand g20 (n_99, A[3], n_97);
  nand g21 (n_100, B[3], n_97);
  nand g22 (n_102, n_98, n_99, n_100);
  xor g23 (n_101, A[3], B[3]);
  xor g24 (Z[3], n_97, n_101);
  nand g25 (n_103, A[4], B[4]);
  nand g26 (n_104, A[4], n_102);
  nand g27 (n_105, B[4], n_102);
  nand g28 (n_107, n_103, n_104, n_105);
  xor g29 (n_106, A[4], B[4]);
  xor g30 (Z[4], n_102, n_106);
  nand g31 (n_108, A[5], B[5]);
  nand g32 (n_109, A[5], n_107);
  nand g33 (n_110, B[5], n_107);
  nand g34 (n_112, n_108, n_109, n_110);
  xor g35 (n_111, A[5], B[5]);
  xor g36 (Z[5], n_107, n_111);
  nand g37 (n_113, A[6], B[6]);
  nand g38 (n_114, A[6], n_112);
  nand g39 (n_115, B[6], n_112);
  nand g40 (n_117, n_113, n_114, n_115);
  xor g41 (n_116, A[6], B[6]);
  xor g42 (Z[6], n_112, n_116);
  nand g43 (n_118, A[7], B[7]);
  nand g44 (n_119, A[7], n_117);
  nand g45 (n_120, B[7], n_117);
  nand g46 (n_122, n_118, n_119, n_120);
  xor g47 (n_121, A[7], B[7]);
  xor g48 (Z[7], n_117, n_121);
  nand g49 (n_123, A[8], B[8]);
  nand g50 (n_124, A[8], n_122);
  nand g51 (n_125, B[8], n_122);
  nand g52 (n_127, n_123, n_124, n_125);
  xor g53 (n_126, A[8], B[8]);
  xor g54 (Z[8], n_122, n_126);
  nand g55 (n_128, A[9], B[9]);
  nand g56 (n_129, A[9], n_127);
  nand g57 (n_130, B[9], n_127);
  nand g58 (n_132, n_128, n_129, n_130);
  xor g59 (n_131, A[9], B[9]);
  xor g60 (Z[9], n_127, n_131);
  nand g61 (n_133, A[10], B[10]);
  nand g62 (n_134, A[10], n_132);
  nand g63 (n_135, B[10], n_132);
  nand g64 (n_137, n_133, n_134, n_135);
  xor g65 (n_136, A[10], B[10]);
  xor g66 (Z[10], n_132, n_136);
  nand g67 (n_138, A[11], B[11]);
  nand g68 (n_139, A[11], n_137);
  nand g69 (n_140, B[11], n_137);
  nand g70 (n_142, n_138, n_139, n_140);
  xor g71 (n_141, A[11], B[11]);
  xor g72 (Z[11], n_137, n_141);
  nand g73 (n_143, A[12], B[12]);
  nand g74 (n_144, A[12], n_142);
  nand g75 (n_145, B[12], n_142);
  nand g76 (n_147, n_143, n_144, n_145);
  xor g77 (n_146, A[12], B[12]);
  xor g78 (Z[12], n_142, n_146);
  nand g79 (n_148, A[13], B[13]);
  nand g80 (n_149, A[13], n_147);
  nand g81 (n_150, B[13], n_147);
  nand g82 (n_152, n_148, n_149, n_150);
  xor g83 (n_151, A[13], B[13]);
  xor g84 (Z[13], n_147, n_151);
  nand g85 (n_153, A[14], B[14]);
  nand g86 (n_154, A[14], n_152);
  nand g87 (n_155, B[14], n_152);
  nand g88 (n_157, n_153, n_154, n_155);
  xor g89 (n_156, A[14], B[14]);
  xor g90 (Z[14], n_152, n_156);
  nand g91 (n_158, A[15], B[15]);
  nand g92 (n_159, A[15], n_157);
  nand g93 (n_160, B[15], n_157);
  nand g94 (n_162, n_158, n_159, n_160);
  xor g95 (n_161, A[15], B[15]);
  xor g96 (Z[15], n_157, n_161);
  nand g97 (n_163, A[16], B[16]);
  nand g98 (n_164, A[16], n_162);
  nand g99 (n_165, B[16], n_162);
  nand g100 (n_167, n_163, n_164, n_165);
  xor g101 (n_166, A[16], B[16]);
  xor g102 (Z[16], n_162, n_166);
  nand g103 (n_168, A[17], B[17]);
  nand g104 (n_169, A[17], n_167);
  nand g105 (n_170, B[17], n_167);
  nand g106 (n_172, n_168, n_169, n_170);
  xor g107 (n_171, A[17], B[17]);
  xor g108 (Z[17], n_167, n_171);
  nand g109 (n_173, A[18], B[18]);
  nand g110 (n_174, A[18], n_172);
  nand g111 (n_175, B[18], n_172);
  nand g112 (n_177, n_173, n_174, n_175);
  xor g113 (n_176, A[18], B[18]);
  xor g114 (Z[18], n_172, n_176);
  nand g115 (n_178, A[19], B[19]);
  nand g116 (n_179, A[19], n_177);
  nand g117 (n_180, B[19], n_177);
  nand g118 (n_182, n_178, n_179, n_180);
  xor g119 (n_181, A[19], B[19]);
  xor g120 (Z[19], n_177, n_181);
  nand g121 (n_183, A[20], B[20]);
  nand g122 (n_184, A[20], n_182);
  nand g123 (n_185, B[20], n_182);
  nand g124 (n_187, n_183, n_184, n_185);
  xor g125 (n_186, A[20], B[20]);
  xor g126 (Z[20], n_182, n_186);
  nand g127 (n_188, A[21], B[21]);
  nand g128 (n_189, A[21], n_187);
  nand g129 (n_190, B[21], n_187);
  nand g130 (n_192, n_188, n_189, n_190);
  xor g131 (n_191, A[21], B[21]);
  xor g132 (Z[21], n_187, n_191);
  nand g133 (n_193, A[22], B[22]);
  nand g134 (n_194, A[22], n_192);
  nand g135 (n_195, B[22], n_192);
  nand g136 (n_197, n_193, n_194, n_195);
  xor g137 (n_196, A[22], B[22]);
  xor g138 (Z[22], n_192, n_196);
  nand g139 (n_198, A[23], B[23]);
  nand g140 (n_199, A[23], n_197);
  nand g141 (n_200, B[23], n_197);
  nand g142 (n_202, n_198, n_199, n_200);
  xor g143 (n_201, A[23], B[23]);
  xor g144 (Z[23], n_197, n_201);
  nand g145 (n_203, A[24], B[24]);
  nand g146 (n_204, A[24], n_202);
  nand g147 (n_205, B[24], n_202);
  nand g148 (n_207, n_203, n_204, n_205);
  xor g149 (n_206, A[24], B[24]);
  xor g150 (Z[24], n_202, n_206);
  nand g151 (n_208, A[25], B[25]);
  nand g152 (n_209, A[25], n_207);
  nand g153 (n_210, B[25], n_207);
  nand g154 (n_212, n_208, n_209, n_210);
  xor g155 (n_211, A[25], B[25]);
  xor g156 (Z[25], n_207, n_211);
  xor g161 (n_216, A[26], B[26]);
  xor g162 (Z[26], n_212, n_216);
  or g164 (n_89, wc, n_83);
  not gc (wc, A[1]);
  or g165 (n_90, wc0, n_83);
  not gc0 (wc0, B[1]);
  xnor g166 (Z[1], n_83, n_91);
endmodule

module add_unsigned_161_GENERIC(A, B, Z);
  input [26:0] A, B;
  output [26:0] Z;
  wire [26:0] A, B;
  wire [26:0] Z;
  add_unsigned_161_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_unsigned_162_GENERIC_REAL(A, B, Z);
// synthesis_equation add_unsigned
  input [26:0] A, B;
  output [26:0] Z;
  wire [26:0] A, B;
  wire [26:0] Z;
  wire n_83, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190;
  wire n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198;
  wire n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_207, n_208, n_209, n_210, n_211, n_212, n_216;
  nand g1 (n_83, A[0], B[0]);
  xor g5 (Z[0], A[0], B[0]);
  nand g7 (n_88, A[1], B[1]);
  nand g10 (n_92, n_88, n_89, n_90);
  xor g11 (n_91, A[1], B[1]);
  nand g13 (n_93, A[2], B[2]);
  nand g14 (n_94, A[2], n_92);
  nand g15 (n_95, B[2], n_92);
  nand g16 (n_97, n_93, n_94, n_95);
  xor g17 (n_96, A[2], B[2]);
  xor g18 (Z[2], n_92, n_96);
  nand g19 (n_98, A[3], B[3]);
  nand g20 (n_99, A[3], n_97);
  nand g21 (n_100, B[3], n_97);
  nand g22 (n_102, n_98, n_99, n_100);
  xor g23 (n_101, A[3], B[3]);
  xor g24 (Z[3], n_97, n_101);
  nand g25 (n_103, A[4], B[4]);
  nand g26 (n_104, A[4], n_102);
  nand g27 (n_105, B[4], n_102);
  nand g28 (n_107, n_103, n_104, n_105);
  xor g29 (n_106, A[4], B[4]);
  xor g30 (Z[4], n_102, n_106);
  nand g31 (n_108, A[5], B[5]);
  nand g32 (n_109, A[5], n_107);
  nand g33 (n_110, B[5], n_107);
  nand g34 (n_112, n_108, n_109, n_110);
  xor g35 (n_111, A[5], B[5]);
  xor g36 (Z[5], n_107, n_111);
  nand g37 (n_113, A[6], B[6]);
  nand g38 (n_114, A[6], n_112);
  nand g39 (n_115, B[6], n_112);
  nand g40 (n_117, n_113, n_114, n_115);
  xor g41 (n_116, A[6], B[6]);
  xor g42 (Z[6], n_112, n_116);
  nand g43 (n_118, A[7], B[7]);
  nand g44 (n_119, A[7], n_117);
  nand g45 (n_120, B[7], n_117);
  nand g46 (n_122, n_118, n_119, n_120);
  xor g47 (n_121, A[7], B[7]);
  xor g48 (Z[7], n_117, n_121);
  nand g49 (n_123, A[8], B[8]);
  nand g50 (n_124, A[8], n_122);
  nand g51 (n_125, B[8], n_122);
  nand g52 (n_127, n_123, n_124, n_125);
  xor g53 (n_126, A[8], B[8]);
  xor g54 (Z[8], n_122, n_126);
  nand g55 (n_128, A[9], B[9]);
  nand g56 (n_129, A[9], n_127);
  nand g57 (n_130, B[9], n_127);
  nand g58 (n_132, n_128, n_129, n_130);
  xor g59 (n_131, A[9], B[9]);
  xor g60 (Z[9], n_127, n_131);
  nand g61 (n_133, A[10], B[10]);
  nand g62 (n_134, A[10], n_132);
  nand g63 (n_135, B[10], n_132);
  nand g64 (n_137, n_133, n_134, n_135);
  xor g65 (n_136, A[10], B[10]);
  xor g66 (Z[10], n_132, n_136);
  nand g67 (n_138, A[11], B[11]);
  nand g68 (n_139, A[11], n_137);
  nand g69 (n_140, B[11], n_137);
  nand g70 (n_142, n_138, n_139, n_140);
  xor g71 (n_141, A[11], B[11]);
  xor g72 (Z[11], n_137, n_141);
  nand g73 (n_143, A[12], B[12]);
  nand g74 (n_144, A[12], n_142);
  nand g75 (n_145, B[12], n_142);
  nand g76 (n_147, n_143, n_144, n_145);
  xor g77 (n_146, A[12], B[12]);
  xor g78 (Z[12], n_142, n_146);
  nand g79 (n_148, A[13], B[13]);
  nand g80 (n_149, A[13], n_147);
  nand g81 (n_150, B[13], n_147);
  nand g82 (n_152, n_148, n_149, n_150);
  xor g83 (n_151, A[13], B[13]);
  xor g84 (Z[13], n_147, n_151);
  nand g85 (n_153, A[14], B[14]);
  nand g86 (n_154, A[14], n_152);
  nand g87 (n_155, B[14], n_152);
  nand g88 (n_157, n_153, n_154, n_155);
  xor g89 (n_156, A[14], B[14]);
  xor g90 (Z[14], n_152, n_156);
  nand g91 (n_158, A[15], B[15]);
  nand g92 (n_159, A[15], n_157);
  nand g93 (n_160, B[15], n_157);
  nand g94 (n_162, n_158, n_159, n_160);
  xor g95 (n_161, A[15], B[15]);
  xor g96 (Z[15], n_157, n_161);
  nand g97 (n_163, A[16], B[16]);
  nand g98 (n_164, A[16], n_162);
  nand g99 (n_165, B[16], n_162);
  nand g100 (n_167, n_163, n_164, n_165);
  xor g101 (n_166, A[16], B[16]);
  xor g102 (Z[16], n_162, n_166);
  nand g103 (n_168, A[17], B[17]);
  nand g104 (n_169, A[17], n_167);
  nand g105 (n_170, B[17], n_167);
  nand g106 (n_172, n_168, n_169, n_170);
  xor g107 (n_171, A[17], B[17]);
  xor g108 (Z[17], n_167, n_171);
  nand g109 (n_173, A[18], B[18]);
  nand g110 (n_174, A[18], n_172);
  nand g111 (n_175, B[18], n_172);
  nand g112 (n_177, n_173, n_174, n_175);
  xor g113 (n_176, A[18], B[18]);
  xor g114 (Z[18], n_172, n_176);
  nand g115 (n_178, A[19], B[19]);
  nand g116 (n_179, A[19], n_177);
  nand g117 (n_180, B[19], n_177);
  nand g118 (n_182, n_178, n_179, n_180);
  xor g119 (n_181, A[19], B[19]);
  xor g120 (Z[19], n_177, n_181);
  nand g121 (n_183, A[20], B[20]);
  nand g122 (n_184, A[20], n_182);
  nand g123 (n_185, B[20], n_182);
  nand g124 (n_187, n_183, n_184, n_185);
  xor g125 (n_186, A[20], B[20]);
  xor g126 (Z[20], n_182, n_186);
  nand g127 (n_188, A[21], B[21]);
  nand g128 (n_189, A[21], n_187);
  nand g129 (n_190, B[21], n_187);
  nand g130 (n_192, n_188, n_189, n_190);
  xor g131 (n_191, A[21], B[21]);
  xor g132 (Z[21], n_187, n_191);
  nand g133 (n_193, A[22], B[22]);
  nand g134 (n_194, A[22], n_192);
  nand g135 (n_195, B[22], n_192);
  nand g136 (n_197, n_193, n_194, n_195);
  xor g137 (n_196, A[22], B[22]);
  xor g138 (Z[22], n_192, n_196);
  nand g139 (n_198, A[23], B[23]);
  nand g140 (n_199, A[23], n_197);
  nand g141 (n_200, B[23], n_197);
  nand g142 (n_202, n_198, n_199, n_200);
  xor g143 (n_201, A[23], B[23]);
  xor g144 (Z[23], n_197, n_201);
  nand g145 (n_203, A[24], B[24]);
  nand g146 (n_204, A[24], n_202);
  nand g147 (n_205, B[24], n_202);
  nand g148 (n_207, n_203, n_204, n_205);
  xor g149 (n_206, A[24], B[24]);
  xor g150 (Z[24], n_202, n_206);
  nand g151 (n_208, A[25], B[25]);
  nand g152 (n_209, A[25], n_207);
  nand g153 (n_210, B[25], n_207);
  nand g154 (n_212, n_208, n_209, n_210);
  xor g155 (n_211, A[25], B[25]);
  xor g156 (Z[25], n_207, n_211);
  xor g161 (n_216, A[26], B[26]);
  xor g162 (Z[26], n_212, n_216);
  or g164 (n_89, wc, n_83);
  not gc (wc, A[1]);
  or g165 (n_90, wc0, n_83);
  not gc0 (wc0, B[1]);
  xnor g166 (Z[1], n_83, n_91);
endmodule

module add_unsigned_162_GENERIC(A, B, Z);
  input [26:0] A, B;
  output [26:0] Z;
  wire [26:0] A, B;
  wire [26:0] Z;
  add_unsigned_162_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_unsigned_carry_358_2_GENERIC_REAL(A, B, CI, Z);
// synthesis_equation add_unsigned_carry
  input [22:0] A, B;
  input CI;
  output [22:0] Z;
  wire [22:0] A, B;
  wire CI;
  wire [22:0] Z;
  wire n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78;
  wire n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86;
  wire n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_184;
  nand g1 (n_71, A[0], B[0]);
  nand g2 (n_72, A[0], CI);
  nand g3 (n_73, B[0], CI);
  nand g4 (n_75, n_71, n_72, n_73);
  xor g5 (n_74, A[0], B[0]);
  xor g6 (Z[0], CI, n_74);
  nand g7 (n_76, A[1], B[1]);
  nand g8 (n_77, A[1], n_75);
  nand g9 (n_78, B[1], n_75);
  nand g10 (n_80, n_76, n_77, n_78);
  xor g11 (n_79, A[1], B[1]);
  xor g12 (Z[1], n_75, n_79);
  nand g13 (n_81, A[2], B[2]);
  nand g14 (n_82, A[2], n_80);
  nand g15 (n_83, B[2], n_80);
  nand g16 (n_85, n_81, n_82, n_83);
  xor g17 (n_84, A[2], B[2]);
  xor g18 (Z[2], n_80, n_84);
  nand g19 (n_86, A[3], B[3]);
  nand g20 (n_87, A[3], n_85);
  nand g21 (n_88, B[3], n_85);
  nand g22 (n_90, n_86, n_87, n_88);
  xor g23 (n_89, A[3], B[3]);
  xor g24 (Z[3], n_85, n_89);
  nand g25 (n_91, A[4], B[4]);
  nand g26 (n_92, A[4], n_90);
  nand g27 (n_93, B[4], n_90);
  nand g28 (n_95, n_91, n_92, n_93);
  xor g29 (n_94, A[4], B[4]);
  xor g30 (Z[4], n_90, n_94);
  nand g31 (n_96, A[5], B[5]);
  nand g32 (n_97, A[5], n_95);
  nand g33 (n_98, B[5], n_95);
  nand g34 (n_100, n_96, n_97, n_98);
  xor g35 (n_99, A[5], B[5]);
  xor g36 (Z[5], n_95, n_99);
  nand g37 (n_101, A[6], B[6]);
  nand g38 (n_102, A[6], n_100);
  nand g39 (n_103, B[6], n_100);
  nand g40 (n_105, n_101, n_102, n_103);
  xor g41 (n_104, A[6], B[6]);
  xor g42 (Z[6], n_100, n_104);
  nand g43 (n_106, A[7], B[7]);
  nand g44 (n_107, A[7], n_105);
  nand g45 (n_108, B[7], n_105);
  nand g46 (n_110, n_106, n_107, n_108);
  xor g47 (n_109, A[7], B[7]);
  xor g48 (Z[7], n_105, n_109);
  nand g49 (n_111, A[8], B[8]);
  nand g50 (n_112, A[8], n_110);
  nand g51 (n_113, B[8], n_110);
  nand g52 (n_115, n_111, n_112, n_113);
  xor g53 (n_114, A[8], B[8]);
  xor g54 (Z[8], n_110, n_114);
  nand g55 (n_116, A[9], B[9]);
  nand g56 (n_117, A[9], n_115);
  nand g57 (n_118, B[9], n_115);
  nand g58 (n_120, n_116, n_117, n_118);
  xor g59 (n_119, A[9], B[9]);
  xor g60 (Z[9], n_115, n_119);
  nand g61 (n_121, A[10], B[10]);
  nand g62 (n_122, A[10], n_120);
  nand g63 (n_123, B[10], n_120);
  nand g64 (n_125, n_121, n_122, n_123);
  xor g65 (n_124, A[10], B[10]);
  xor g66 (Z[10], n_120, n_124);
  nand g67 (n_126, A[11], B[11]);
  nand g68 (n_127, A[11], n_125);
  nand g69 (n_128, B[11], n_125);
  nand g70 (n_130, n_126, n_127, n_128);
  xor g71 (n_129, A[11], B[11]);
  xor g72 (Z[11], n_125, n_129);
  nand g73 (n_131, A[12], B[12]);
  nand g74 (n_132, A[12], n_130);
  nand g75 (n_133, B[12], n_130);
  nand g76 (n_135, n_131, n_132, n_133);
  xor g77 (n_134, A[12], B[12]);
  xor g78 (Z[12], n_130, n_134);
  nand g79 (n_136, A[13], B[13]);
  nand g80 (n_137, A[13], n_135);
  nand g81 (n_138, B[13], n_135);
  nand g82 (n_140, n_136, n_137, n_138);
  xor g83 (n_139, A[13], B[13]);
  xor g84 (Z[13], n_135, n_139);
  nand g85 (n_141, A[14], B[14]);
  nand g86 (n_142, A[14], n_140);
  nand g87 (n_143, B[14], n_140);
  nand g88 (n_145, n_141, n_142, n_143);
  xor g89 (n_144, A[14], B[14]);
  xor g90 (Z[14], n_140, n_144);
  nand g91 (n_146, A[15], B[15]);
  nand g92 (n_147, A[15], n_145);
  nand g93 (n_148, B[15], n_145);
  nand g94 (n_150, n_146, n_147, n_148);
  xor g95 (n_149, A[15], B[15]);
  xor g96 (Z[15], n_145, n_149);
  nand g97 (n_151, A[16], B[16]);
  nand g98 (n_152, A[16], n_150);
  nand g99 (n_153, B[16], n_150);
  nand g100 (n_155, n_151, n_152, n_153);
  xor g101 (n_154, A[16], B[16]);
  xor g102 (Z[16], n_150, n_154);
  nand g103 (n_156, A[17], B[17]);
  nand g104 (n_157, A[17], n_155);
  nand g105 (n_158, B[17], n_155);
  nand g106 (n_160, n_156, n_157, n_158);
  xor g107 (n_159, A[17], B[17]);
  xor g108 (Z[17], n_155, n_159);
  nand g109 (n_161, A[18], B[18]);
  nand g110 (n_162, A[18], n_160);
  nand g111 (n_163, B[18], n_160);
  nand g112 (n_165, n_161, n_162, n_163);
  xor g113 (n_164, A[18], B[18]);
  xor g114 (Z[18], n_160, n_164);
  nand g115 (n_166, A[19], B[19]);
  nand g116 (n_167, A[19], n_165);
  nand g117 (n_168, B[19], n_165);
  nand g118 (n_170, n_166, n_167, n_168);
  xor g119 (n_169, A[19], B[19]);
  xor g120 (Z[19], n_165, n_169);
  nand g121 (n_171, A[20], B[20]);
  nand g122 (n_172, A[20], n_170);
  nand g123 (n_173, B[20], n_170);
  nand g124 (n_175, n_171, n_172, n_173);
  xor g125 (n_174, A[20], B[20]);
  xor g126 (Z[20], n_170, n_174);
  nand g127 (n_176, A[21], B[21]);
  nand g128 (n_177, A[21], n_175);
  nand g129 (n_178, B[21], n_175);
  nand g130 (n_180, n_176, n_177, n_178);
  xor g131 (n_179, A[21], B[21]);
  xor g132 (Z[21], n_175, n_179);
  xor g137 (n_184, A[22], B[22]);
  xor g138 (Z[22], n_180, n_184);
endmodule

module add_unsigned_carry_358_2_GENERIC(A, B, CI, Z);
  input [22:0] A, B;
  input CI;
  output [22:0] Z;
  wire [22:0] A, B;
  wire CI;
  wire [22:0] Z;
  wire n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8;
  wire n_9, n_10, n_11, n_12, n_13, n_14, n_15, n_16;
  wire n_17, n_18, n_19, n_20, n_21, n_45;
  add_unsigned_carry_358_2_GENERIC_REAL g1(.A ({n_1, n_2, n_3, n_4,
       n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15,
       n_16, n_17, n_18, n_19, n_20, n_21, A[1:0]}), .B ({B[22:2],
       n_45, B[0]}), .CI (CI), .Z (Z));
  not g2 (n_1, B[21]);
  not g3 (n_2, B[20]);
  not g4 (n_3, B[19]);
  not g5 (n_4, B[18]);
  not g6 (n_5, B[17]);
  not g7 (n_6, B[16]);
  not g8 (n_7, B[15]);
  not g9 (n_8, B[14]);
  not g10 (n_9, B[13]);
  not g11 (n_10, B[12]);
  not g12 (n_11, B[11]);
  not g13 (n_12, B[10]);
  not g14 (n_13, B[9]);
  not g15 (n_14, B[8]);
  not g16 (n_15, B[7]);
  not g17 (n_16, B[6]);
  not g18 (n_17, B[5]);
  not g19 (n_18, B[4]);
  not g20 (n_19, B[3]);
  not g21 (n_20, B[2]);
  not g22 (n_21, A[1]);
  not g23 (n_45, B[0]);
endmodule

module csa_tree_308_GENERIC_REAL(in_0, out_0, out_1);
// synthesis_equation "assign out_0 = ( $signed({1'b0,in_0}) - 128 )  ; assign out_1 = 10'b0;"
  input [7:0] in_0;
  output [9:0] out_0, out_1;
  wire [7:0] in_0;
  wire [9:0] out_0, out_1;
  assign out_1[0] = 1'b0;
  assign out_1[1] = 1'b0;
  assign out_1[2] = 1'b0;
  assign out_1[3] = 1'b0;
  assign out_1[4] = 1'b0;
  assign out_1[5] = 1'b0;
  assign out_1[6] = 1'b0;
  assign out_1[7] = 1'b1;
  assign out_1[8] = 1'b0;
  assign out_1[9] = 1'b0;
  assign out_0[0] = in_0[0];
  assign out_0[1] = in_0[1];
  assign out_0[2] = in_0[2];
  assign out_0[3] = in_0[3];
  assign out_0[4] = in_0[4];
  assign out_0[5] = in_0[5];
  assign out_0[6] = in_0[6];
  assign out_0[7] = in_0[7];
  assign out_0[8] = 1'b1;
  assign out_0[9] = 1'b1;
endmodule

module csa_tree_308_GENERIC(in_0, out_0, out_1);
  input [7:0] in_0;
  output [9:0] out_0, out_1;
  wire [7:0] in_0;
  wire [9:0] out_0, out_1;
  csa_tree_308_GENERIC_REAL g1(.in_0 (in_0), .out_0 (out_0), .out_1
       (out_1));
endmodule

module csa_tree_308_1_GENERIC_REAL(in_0, out_0, out_1);
// synthesis_equation "assign out_0 = ( $signed({1'b0,in_0}) - 128 )  ; assign out_1 = 10'b0;"
  input [7:0] in_0;
  output [9:0] out_0, out_1;
  wire [7:0] in_0;
  wire [9:0] out_0, out_1;
  assign out_1[0] = 1'b0;
  assign out_1[1] = 1'b0;
  assign out_1[2] = 1'b0;
  assign out_1[3] = 1'b0;
  assign out_1[4] = 1'b0;
  assign out_1[5] = 1'b0;
  assign out_1[6] = 1'b0;
  assign out_1[7] = 1'b1;
  assign out_1[8] = 1'b0;
  assign out_1[9] = 1'b0;
  assign out_0[0] = in_0[0];
  assign out_0[1] = in_0[1];
  assign out_0[2] = in_0[2];
  assign out_0[3] = in_0[3];
  assign out_0[4] = in_0[4];
  assign out_0[5] = in_0[5];
  assign out_0[6] = in_0[6];
  assign out_0[7] = in_0[7];
  assign out_0[8] = 1'b1;
  assign out_0[9] = 1'b1;
endmodule

module csa_tree_308_1_GENERIC(in_0, out_0, out_1);
  input [7:0] in_0;
  output [9:0] out_0, out_1;
  wire [7:0] in_0;
  wire [9:0] out_0, out_1;
  csa_tree_308_1_GENERIC_REAL g1(.in_0 (in_0), .out_0 (out_0), .out_1
       (out_1));
endmodule

module increment_unsigned_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [24:0] A;
  input CI;
  output [24:0] Z;
  wire [24:0] A;
  wire CI;
  wire [24:0] Z;
  wire n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59;
  wire n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67;
  wire n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_52, A[0], CI);
  xor g25 (Z[1], A[1], n_52);
  and g26 (n_53, A[1], n_52);
  xor g27 (Z[2], A[2], n_53);
  and g28 (n_54, A[2], n_53);
  xor g29 (Z[3], A[3], n_54);
  and g30 (n_55, A[3], n_54);
  xor g31 (Z[4], A[4], n_55);
  and g32 (n_56, A[4], n_55);
  xor g33 (Z[5], A[5], n_56);
  and g34 (n_57, A[5], n_56);
  xor g35 (Z[6], A[6], n_57);
  and g36 (n_58, A[6], n_57);
  xor g37 (Z[7], A[7], n_58);
  and g38 (n_59, A[7], n_58);
  xor g39 (Z[8], A[8], n_59);
  and g40 (n_60, A[8], n_59);
  xor g41 (Z[9], A[9], n_60);
  and g42 (n_61, A[9], n_60);
  xor g43 (Z[10], A[10], n_61);
  and g44 (n_62, A[10], n_61);
  xor g45 (Z[11], A[11], n_62);
  and g46 (n_63, A[11], n_62);
  xor g47 (Z[12], A[12], n_63);
  and g48 (n_64, A[12], n_63);
  xor g49 (Z[13], A[13], n_64);
  and g50 (n_65, A[13], n_64);
  xor g51 (Z[14], A[14], n_65);
  and g52 (n_66, A[14], n_65);
  xor g53 (Z[15], A[15], n_66);
  and g54 (n_67, A[15], n_66);
  xor g55 (Z[16], A[16], n_67);
  and g56 (n_68, A[16], n_67);
  xor g57 (Z[17], A[17], n_68);
  and g58 (n_69, A[17], n_68);
  xor g59 (Z[18], A[18], n_69);
  and g60 (n_70, A[18], n_69);
  xor g61 (Z[19], A[19], n_70);
  and g62 (n_71, A[19], n_70);
  xor g63 (Z[20], A[20], n_71);
  and g64 (n_72, A[20], n_71);
  xor g65 (Z[21], A[21], n_72);
  and g66 (n_73, A[21], n_72);
  xor g67 (Z[22], A[22], n_73);
  and g68 (n_74, A[22], n_73);
  xor g69 (Z[23], A[23], n_74);
  and g70 (n_75, A[23], n_74);
  xor g71 (Z[24], A[24], n_75);
endmodule

module increment_unsigned_GENERIC(A, CI, Z);
  input [24:0] A;
  input CI;
  output [24:0] Z;
  wire [24:0] A;
  wire CI;
  wire [24:0] Z;
  increment_unsigned_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_1_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [24:0] A;
  input CI;
  output [24:0] Z;
  wire [24:0] A;
  wire CI;
  wire [24:0] Z;
  wire n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59;
  wire n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67;
  wire n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_52, A[0], CI);
  xor g25 (Z[1], A[1], n_52);
  and g26 (n_53, A[1], n_52);
  xor g27 (Z[2], A[2], n_53);
  and g28 (n_54, A[2], n_53);
  xor g29 (Z[3], A[3], n_54);
  and g30 (n_55, A[3], n_54);
  xor g31 (Z[4], A[4], n_55);
  and g32 (n_56, A[4], n_55);
  xor g33 (Z[5], A[5], n_56);
  and g34 (n_57, A[5], n_56);
  xor g35 (Z[6], A[6], n_57);
  and g36 (n_58, A[6], n_57);
  xor g37 (Z[7], A[7], n_58);
  and g38 (n_59, A[7], n_58);
  xor g39 (Z[8], A[8], n_59);
  and g40 (n_60, A[8], n_59);
  xor g41 (Z[9], A[9], n_60);
  and g42 (n_61, A[9], n_60);
  xor g43 (Z[10], A[10], n_61);
  and g44 (n_62, A[10], n_61);
  xor g45 (Z[11], A[11], n_62);
  and g46 (n_63, A[11], n_62);
  xor g47 (Z[12], A[12], n_63);
  and g48 (n_64, A[12], n_63);
  xor g49 (Z[13], A[13], n_64);
  and g50 (n_65, A[13], n_64);
  xor g51 (Z[14], A[14], n_65);
  and g52 (n_66, A[14], n_65);
  xor g53 (Z[15], A[15], n_66);
  and g54 (n_67, A[15], n_66);
  xor g55 (Z[16], A[16], n_67);
  and g56 (n_68, A[16], n_67);
  xor g57 (Z[17], A[17], n_68);
  and g58 (n_69, A[17], n_68);
  xor g59 (Z[18], A[18], n_69);
  and g60 (n_70, A[18], n_69);
  xor g61 (Z[19], A[19], n_70);
  and g62 (n_71, A[19], n_70);
  xor g63 (Z[20], A[20], n_71);
  and g64 (n_72, A[20], n_71);
  xor g65 (Z[21], A[21], n_72);
  and g66 (n_73, A[21], n_72);
  xor g67 (Z[22], A[22], n_73);
  and g68 (n_74, A[22], n_73);
  xor g69 (Z[23], A[23], n_74);
  and g70 (n_75, A[23], n_74);
  xor g71 (Z[24], A[24], n_75);
endmodule

module increment_unsigned_1_GENERIC(A, CI, Z);
  input [24:0] A;
  input CI;
  output [24:0] Z;
  wire [24:0] A;
  wire CI;
  wire [24:0] Z;
  increment_unsigned_1_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_1_1252_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [24:0] A;
  input CI;
  output [24:0] Z;
  wire [24:0] A;
  wire CI;
  wire [24:0] Z;
  wire n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59;
  wire n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67;
  wire n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_52, A[0], CI);
  xor g25 (Z[1], A[1], n_52);
  and g26 (n_53, A[1], n_52);
  xor g27 (Z[2], A[2], n_53);
  and g28 (n_54, A[2], n_53);
  xor g29 (Z[3], A[3], n_54);
  and g30 (n_55, A[3], n_54);
  xor g31 (Z[4], A[4], n_55);
  and g32 (n_56, A[4], n_55);
  xor g33 (Z[5], A[5], n_56);
  and g34 (n_57, A[5], n_56);
  xor g35 (Z[6], A[6], n_57);
  and g36 (n_58, A[6], n_57);
  xor g37 (Z[7], A[7], n_58);
  and g38 (n_59, A[7], n_58);
  xor g39 (Z[8], A[8], n_59);
  and g40 (n_60, A[8], n_59);
  xor g41 (Z[9], A[9], n_60);
  and g42 (n_61, A[9], n_60);
  xor g43 (Z[10], A[10], n_61);
  and g44 (n_62, A[10], n_61);
  xor g45 (Z[11], A[11], n_62);
  and g46 (n_63, A[11], n_62);
  xor g47 (Z[12], A[12], n_63);
  and g48 (n_64, A[12], n_63);
  xor g49 (Z[13], A[13], n_64);
  and g50 (n_65, A[13], n_64);
  xor g51 (Z[14], A[14], n_65);
  and g52 (n_66, A[14], n_65);
  xor g53 (Z[15], A[15], n_66);
  and g54 (n_67, A[15], n_66);
  xor g55 (Z[16], A[16], n_67);
  and g56 (n_68, A[16], n_67);
  xor g57 (Z[17], A[17], n_68);
  and g58 (n_69, A[17], n_68);
  xor g59 (Z[18], A[18], n_69);
  and g60 (n_70, A[18], n_69);
  xor g61 (Z[19], A[19], n_70);
  and g62 (n_71, A[19], n_70);
  xor g63 (Z[20], A[20], n_71);
  and g64 (n_72, A[20], n_71);
  xor g65 (Z[21], A[21], n_72);
  and g66 (n_73, A[21], n_72);
  xor g67 (Z[22], A[22], n_73);
  and g68 (n_74, A[22], n_73);
  xor g69 (Z[23], A[23], n_74);
  and g70 (n_75, A[23], n_74);
  xor g71 (Z[24], A[24], n_75);
endmodule

module increment_unsigned_1_1252_GENERIC(A, CI, Z);
  input [24:0] A;
  input CI;
  output [24:0] Z;
  wire [24:0] A;
  wire CI;
  wire [24:0] Z;
  increment_unsigned_1_1252_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_332_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [26:0] A;
  input CI;
  output [26:0] Z;
  wire [26:0] A;
  wire CI;
  wire [26:0] Z;
  wire n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63;
  wire n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71;
  wire n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79;
  wire n_80, n_81;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_56, A[0], CI);
  xor g27 (Z[1], A[1], n_56);
  and g28 (n_57, A[1], n_56);
  xor g29 (Z[2], A[2], n_57);
  and g30 (n_58, A[2], n_57);
  xor g31 (Z[3], A[3], n_58);
  and g32 (n_59, A[3], n_58);
  xor g33 (Z[4], A[4], n_59);
  and g34 (n_60, A[4], n_59);
  xor g35 (Z[5], A[5], n_60);
  and g36 (n_61, A[5], n_60);
  xor g37 (Z[6], A[6], n_61);
  and g38 (n_62, A[6], n_61);
  xor g39 (Z[7], A[7], n_62);
  and g40 (n_63, A[7], n_62);
  xor g41 (Z[8], A[8], n_63);
  and g42 (n_64, A[8], n_63);
  xor g43 (Z[9], A[9], n_64);
  and g44 (n_65, A[9], n_64);
  xor g45 (Z[10], A[10], n_65);
  and g46 (n_66, A[10], n_65);
  xor g47 (Z[11], A[11], n_66);
  and g48 (n_67, A[11], n_66);
  xor g49 (Z[12], A[12], n_67);
  and g50 (n_68, A[12], n_67);
  xor g51 (Z[13], A[13], n_68);
  and g52 (n_69, A[13], n_68);
  xor g53 (Z[14], A[14], n_69);
  and g54 (n_70, A[14], n_69);
  xor g55 (Z[15], A[15], n_70);
  and g56 (n_71, A[15], n_70);
  xor g57 (Z[16], A[16], n_71);
  and g58 (n_72, A[16], n_71);
  xor g59 (Z[17], A[17], n_72);
  and g60 (n_73, A[17], n_72);
  xor g61 (Z[18], A[18], n_73);
  and g62 (n_74, A[18], n_73);
  xor g63 (Z[19], A[19], n_74);
  and g64 (n_75, A[19], n_74);
  xor g65 (Z[20], A[20], n_75);
  and g66 (n_76, A[20], n_75);
  xor g67 (Z[21], A[21], n_76);
  and g68 (n_77, A[21], n_76);
  xor g69 (Z[22], A[22], n_77);
  and g70 (n_78, A[22], n_77);
  xor g71 (Z[23], A[23], n_78);
  and g72 (n_79, A[23], n_78);
  xor g73 (Z[24], A[24], n_79);
  and g74 (n_80, A[24], n_79);
  xor g75 (Z[25], A[25], n_80);
  and g76 (n_81, A[25], n_80);
  xor g77 (Z[26], A[26], n_81);
endmodule

module increment_unsigned_332_GENERIC(A, CI, Z);
  input [26:0] A;
  input CI;
  output [26:0] Z;
  wire [26:0] A;
  wire CI;
  wire [26:0] Z;
  increment_unsigned_332_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_355_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [22:0] A;
  input CI;
  output [22:0] Z;
  wire [22:0] A;
  wire CI;
  wire [22:0] Z;
  wire n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55;
  wire n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63;
  wire n_64, n_65, n_66, n_67, n_68, n_69;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_48, A[0], CI);
  xor g23 (Z[1], A[1], n_48);
  and g24 (n_49, A[1], n_48);
  xor g25 (Z[2], A[2], n_49);
  and g26 (n_50, A[2], n_49);
  xor g27 (Z[3], A[3], n_50);
  and g28 (n_51, A[3], n_50);
  xor g29 (Z[4], A[4], n_51);
  and g30 (n_52, A[4], n_51);
  xor g31 (Z[5], A[5], n_52);
  and g32 (n_53, A[5], n_52);
  xor g33 (Z[6], A[6], n_53);
  and g34 (n_54, A[6], n_53);
  xor g35 (Z[7], A[7], n_54);
  and g36 (n_55, A[7], n_54);
  xor g37 (Z[8], A[8], n_55);
  and g38 (n_56, A[8], n_55);
  xor g39 (Z[9], A[9], n_56);
  and g40 (n_57, A[9], n_56);
  xor g41 (Z[10], A[10], n_57);
  and g42 (n_58, A[10], n_57);
  xor g43 (Z[11], A[11], n_58);
  and g44 (n_59, A[11], n_58);
  xor g45 (Z[12], A[12], n_59);
  and g46 (n_60, A[12], n_59);
  xor g47 (Z[13], A[13], n_60);
  and g48 (n_61, A[13], n_60);
  xor g49 (Z[14], A[14], n_61);
  and g50 (n_62, A[14], n_61);
  xor g51 (Z[15], A[15], n_62);
  and g52 (n_63, A[15], n_62);
  xor g53 (Z[16], A[16], n_63);
  and g54 (n_64, A[16], n_63);
  xor g55 (Z[17], A[17], n_64);
  and g56 (n_65, A[17], n_64);
  xor g57 (Z[18], A[18], n_65);
  and g58 (n_66, A[18], n_65);
  xor g59 (Z[19], A[19], n_66);
  and g60 (n_67, A[19], n_66);
  xor g61 (Z[20], A[20], n_67);
  and g62 (n_68, A[20], n_67);
  xor g63 (Z[21], A[21], n_68);
  and g64 (n_69, A[21], n_68);
  xor g65 (Z[22], A[22], n_69);
endmodule

module increment_unsigned_355_GENERIC(A, CI, Z);
  input [22:0] A;
  input CI;
  output [22:0] Z;
  wire [22:0] A;
  wire CI;
  wire [22:0] Z;
  increment_unsigned_355_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_355_1_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [22:0] A;
  input CI;
  output [22:0] Z;
  wire [22:0] A;
  wire CI;
  wire [22:0] Z;
  wire n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55;
  wire n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63;
  wire n_64, n_65, n_66, n_67, n_68, n_69;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_48, A[0], CI);
  xor g23 (Z[1], A[1], n_48);
  and g24 (n_49, A[1], n_48);
  xor g25 (Z[2], A[2], n_49);
  and g26 (n_50, A[2], n_49);
  xor g27 (Z[3], A[3], n_50);
  and g28 (n_51, A[3], n_50);
  xor g29 (Z[4], A[4], n_51);
  and g30 (n_52, A[4], n_51);
  xor g31 (Z[5], A[5], n_52);
  and g32 (n_53, A[5], n_52);
  xor g33 (Z[6], A[6], n_53);
  and g34 (n_54, A[6], n_53);
  xor g35 (Z[7], A[7], n_54);
  and g36 (n_55, A[7], n_54);
  xor g37 (Z[8], A[8], n_55);
  and g38 (n_56, A[8], n_55);
  xor g39 (Z[9], A[9], n_56);
  and g40 (n_57, A[9], n_56);
  xor g41 (Z[10], A[10], n_57);
  and g42 (n_58, A[10], n_57);
  xor g43 (Z[11], A[11], n_58);
  and g44 (n_59, A[11], n_58);
  xor g45 (Z[12], A[12], n_59);
  and g46 (n_60, A[12], n_59);
  xor g47 (Z[13], A[13], n_60);
  and g48 (n_61, A[13], n_60);
  xor g49 (Z[14], A[14], n_61);
  and g50 (n_62, A[14], n_61);
  xor g51 (Z[15], A[15], n_62);
  and g52 (n_63, A[15], n_62);
  xor g53 (Z[16], A[16], n_63);
  and g54 (n_64, A[16], n_63);
  xor g55 (Z[17], A[17], n_64);
  and g56 (n_65, A[17], n_64);
  xor g57 (Z[18], A[18], n_65);
  and g58 (n_66, A[18], n_65);
  xor g59 (Z[19], A[19], n_66);
  and g60 (n_67, A[19], n_66);
  xor g61 (Z[20], A[20], n_67);
  and g62 (n_68, A[20], n_67);
  xor g63 (Z[21], A[21], n_68);
  and g64 (n_69, A[21], n_68);
  xor g65 (Z[22], A[22], n_69);
endmodule

module increment_unsigned_355_1_GENERIC(A, CI, Z);
  input [22:0] A;
  input CI;
  output [22:0] Z;
  wire [22:0] A;
  wire CI;
  wire [22:0] Z;
  increment_unsigned_355_1_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_355_2_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [22:0] A;
  input CI;
  output [22:0] Z;
  wire [22:0] A;
  wire CI;
  wire [22:0] Z;
  wire n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55;
  wire n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63;
  wire n_64, n_65, n_66, n_67, n_68, n_69;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_48, A[0], CI);
  xor g23 (Z[1], A[1], n_48);
  and g24 (n_49, A[1], n_48);
  xor g25 (Z[2], A[2], n_49);
  and g26 (n_50, A[2], n_49);
  xor g27 (Z[3], A[3], n_50);
  and g28 (n_51, A[3], n_50);
  xor g29 (Z[4], A[4], n_51);
  and g30 (n_52, A[4], n_51);
  xor g31 (Z[5], A[5], n_52);
  and g32 (n_53, A[5], n_52);
  xor g33 (Z[6], A[6], n_53);
  and g34 (n_54, A[6], n_53);
  xor g35 (Z[7], A[7], n_54);
  and g36 (n_55, A[7], n_54);
  xor g37 (Z[8], A[8], n_55);
  and g38 (n_56, A[8], n_55);
  xor g39 (Z[9], A[9], n_56);
  and g40 (n_57, A[9], n_56);
  xor g41 (Z[10], A[10], n_57);
  and g42 (n_58, A[10], n_57);
  xor g43 (Z[11], A[11], n_58);
  and g44 (n_59, A[11], n_58);
  xor g45 (Z[12], A[12], n_59);
  and g46 (n_60, A[12], n_59);
  xor g47 (Z[13], A[13], n_60);
  and g48 (n_61, A[13], n_60);
  xor g49 (Z[14], A[14], n_61);
  and g50 (n_62, A[14], n_61);
  xor g51 (Z[15], A[15], n_62);
  and g52 (n_63, A[15], n_62);
  xor g53 (Z[16], A[16], n_63);
  and g54 (n_64, A[16], n_63);
  xor g55 (Z[17], A[17], n_64);
  and g56 (n_65, A[17], n_64);
  xor g57 (Z[18], A[18], n_65);
  and g58 (n_66, A[18], n_65);
  xor g59 (Z[19], A[19], n_66);
  and g60 (n_67, A[19], n_66);
  xor g61 (Z[20], A[20], n_67);
  and g62 (n_68, A[20], n_67);
  xor g63 (Z[21], A[21], n_68);
  and g64 (n_69, A[21], n_68);
  xor g65 (Z[22], A[22], n_69);
endmodule

module increment_unsigned_355_2_GENERIC(A, CI, Z);
  input [22:0] A;
  input CI;
  output [22:0] Z;
  wire [22:0] A;
  wire CI;
  wire [22:0] Z;
  increment_unsigned_355_2_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module mult_unsigned_GENERIC_REAL(A, B, Z);
// synthesis_equation "assign Z = $unsigned(A) * $unsigned(B);"
  input [25:0] A, B;
  output [51:0] Z;
  wire [25:0] A, B;
  wire [51:0] Z;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_197, n_198, n_199, n_200, n_201, n_202, n_204, n_311;
  wire n_313, n_315, n_319, n_322, n_323, n_324, n_325, n_326;
  wire n_327, n_328, n_329, n_330, n_331, n_332, n_333, n_334;
  wire n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342;
  wire n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350;
  wire n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366;
  wire n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_391, n_392, n_393, n_396, n_397, n_401, n_402, n_404;
  wire n_405, n_406, n_407, n_408, n_410, n_412, n_416, n_419;
  wire n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427;
  wire n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435;
  wire n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443;
  wire n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451;
  wire n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459;
  wire n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467;
  wire n_468, n_469, n_470, n_471, n_472, n_473, n_474, n_475;
  wire n_476, n_477, n_478, n_479, n_480, n_481, n_482, n_483;
  wire n_484, n_485, n_486, n_487, n_488, n_489, n_490, n_493;
  wire n_494, n_498, n_499, n_501, n_502, n_503, n_504, n_505;
  wire n_507, n_509, n_513, n_516, n_517, n_518, n_519, n_520;
  wire n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528;
  wire n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536;
  wire n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544;
  wire n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552;
  wire n_553, n_554, n_555, n_556, n_557, n_558, n_559, n_560;
  wire n_561, n_562, n_563, n_564, n_565, n_566, n_567, n_568;
  wire n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576;
  wire n_577, n_578, n_579, n_580, n_581, n_582, n_583, n_584;
  wire n_585, n_586, n_587, n_590, n_591, n_595, n_596, n_598;
  wire n_599, n_600, n_601, n_602, n_604, n_606, n_610, n_613;
  wire n_614, n_615, n_616, n_617, n_618, n_619, n_620, n_621;
  wire n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629;
  wire n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637;
  wire n_638, n_639, n_640, n_641, n_642, n_643, n_644, n_645;
  wire n_646, n_647, n_648, n_649, n_650, n_651, n_652, n_653;
  wire n_654, n_655, n_656, n_657, n_658, n_659, n_660, n_661;
  wire n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_669;
  wire n_670, n_671, n_672, n_673, n_674, n_675, n_676, n_677;
  wire n_678, n_679, n_680, n_681, n_682, n_683, n_684, n_687;
  wire n_688, n_692, n_693, n_695, n_696, n_697, n_698, n_699;
  wire n_701, n_703, n_707, n_710, n_711, n_712, n_713, n_714;
  wire n_715, n_716, n_717, n_718, n_719, n_720, n_721, n_722;
  wire n_723, n_724, n_725, n_726, n_727, n_728, n_729, n_730;
  wire n_731, n_732, n_733, n_734, n_735, n_736, n_737, n_738;
  wire n_739, n_740, n_741, n_742, n_743, n_744, n_745, n_746;
  wire n_747, n_748, n_749, n_750, n_751, n_752, n_753, n_754;
  wire n_755, n_756, n_757, n_758, n_759, n_760, n_761, n_762;
  wire n_763, n_764, n_765, n_766, n_767, n_768, n_769, n_770;
  wire n_771, n_772, n_773, n_774, n_775, n_776, n_777, n_778;
  wire n_779, n_780, n_781, n_784, n_785, n_789, n_790, n_792;
  wire n_793, n_794, n_795, n_796, n_798, n_800, n_804, n_807;
  wire n_808, n_809, n_810, n_811, n_812, n_813, n_814, n_815;
  wire n_816, n_817, n_818, n_819, n_820, n_821, n_822, n_823;
  wire n_824, n_825, n_826, n_827, n_828, n_829, n_830, n_831;
  wire n_832, n_833, n_834, n_835, n_836, n_837, n_838, n_839;
  wire n_840, n_841, n_842, n_843, n_844, n_845, n_846, n_847;
  wire n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855;
  wire n_856, n_857, n_858, n_859, n_860, n_861, n_862, n_863;
  wire n_864, n_865, n_866, n_867, n_868, n_869, n_870, n_871;
  wire n_872, n_873, n_874, n_875, n_876, n_877, n_878, n_881;
  wire n_882, n_886, n_887, n_889, n_890, n_891, n_892, n_893;
  wire n_895, n_897, n_901, n_904, n_905, n_906, n_907, n_908;
  wire n_909, n_910, n_911, n_912, n_913, n_914, n_915, n_916;
  wire n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924;
  wire n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932;
  wire n_933, n_934, n_935, n_936, n_937, n_938, n_939, n_940;
  wire n_941, n_942, n_943, n_944, n_945, n_946, n_947, n_948;
  wire n_949, n_950, n_951, n_952, n_953, n_954, n_955, n_956;
  wire n_957, n_958, n_959, n_960, n_961, n_962, n_963, n_964;
  wire n_965, n_966, n_967, n_968, n_969, n_970, n_971, n_972;
  wire n_973, n_974, n_975, n_978, n_979, n_983, n_984, n_986;
  wire n_987, n_988, n_989, n_990, n_992, n_994, n_998, n_1001;
  wire n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009;
  wire n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017;
  wire n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025;
  wire n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033;
  wire n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041;
  wire n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049;
  wire n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057;
  wire n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065;
  wire n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1075;
  wire n_1076, n_1080, n_1081, n_1083, n_1084, n_1085, n_1086, n_1087;
  wire n_1089, n_1091, n_1095, n_1098, n_1099, n_1100, n_1101, n_1102;
  wire n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110;
  wire n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118;
  wire n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126;
  wire n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134;
  wire n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142;
  wire n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150;
  wire n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158;
  wire n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166;
  wire n_1167, n_1168, n_1169, n_1172, n_1173, n_1177, n_1178, n_1180;
  wire n_1181, n_1182, n_1183, n_1184, n_1186, n_1188, n_1192, n_1195;
  wire n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203;
  wire n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211;
  wire n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219;
  wire n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227;
  wire n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235;
  wire n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243;
  wire n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251;
  wire n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259;
  wire n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1269;
  wire n_1270, n_1274, n_1275, n_1277, n_1278, n_1279, n_1280, n_1281;
  wire n_1283, n_1285, n_1289, n_1292, n_1293, n_1294, n_1295, n_1296;
  wire n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304;
  wire n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312;
  wire n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320;
  wire n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328;
  wire n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336;
  wire n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344;
  wire n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352;
  wire n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360;
  wire n_1361, n_1362, n_1363, n_1366, n_1367, n_1371, n_1372, n_1374;
  wire n_1375, n_1376, n_1377, n_1378, n_1380, n_1382, n_1386, n_1389;
  wire n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397;
  wire n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405;
  wire n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413;
  wire n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421;
  wire n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429;
  wire n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437;
  wire n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445;
  wire n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453;
  wire n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1463;
  wire n_1464, n_1468, n_1469, n_1471, n_1472, n_1473, n_1474, n_1497;
  wire n_1501, n_1505, n_1509, n_1513, n_1517, n_1521, n_1525, n_1529;
  wire n_1533, n_1537, n_1541, n_1545, n_1549, n_1553, n_1557, n_1561;
  wire n_1565, n_1569, n_1573, n_1577, n_1581, n_1585, n_1597, n_1598;
  wire n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606;
  wire n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614;
  wire n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622;
  wire n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630;
  wire n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638;
  wire n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646;
  wire n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654;
  wire n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662;
  wire n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670;
  wire n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678;
  wire n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686;
  wire n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694;
  wire n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702;
  wire n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710;
  wire n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718;
  wire n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726;
  wire n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734;
  wire n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742;
  wire n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750;
  wire n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758;
  wire n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766;
  wire n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774;
  wire n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782;
  wire n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790;
  wire n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798;
  wire n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806;
  wire n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814;
  wire n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822;
  wire n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830;
  wire n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838;
  wire n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846;
  wire n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854;
  wire n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862;
  wire n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870;
  wire n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878;
  wire n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886;
  wire n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894;
  wire n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902;
  wire n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910;
  wire n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918;
  wire n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926;
  wire n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934;
  wire n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942;
  wire n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950;
  wire n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958;
  wire n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966;
  wire n_1967, n_1968, n_1969, n_1970, n_1972, n_1973, n_1974, n_1975;
  wire n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983;
  wire n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991;
  wire n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999;
  wire n_2000, n_2001, n_2002, n_2003, n_2006, n_2007, n_2008, n_2009;
  wire n_2010, n_2011, n_2013, n_2014, n_2015, n_2016, n_2017, n_2019;
  wire n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027;
  wire n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035;
  wire n_2036, n_2037, n_2038, n_2041, n_2042, n_2043, n_2044, n_2045;
  wire n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2054, n_2055;
  wire n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063;
  wire n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071;
  wire n_2072, n_2073, n_2075, n_2076, n_2078, n_2079, n_2080, n_2081;
  wire n_2082, n_2083, n_2084, n_2085, n_2087, n_2088, n_2089, n_2090;
  wire n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098;
  wire n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106;
  wire n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116;
  wire n_2117, n_2118, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125;
  wire n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133;
  wire n_2134, n_2135, n_2136, n_2137, n_2138, n_2140, n_2141, n_2143;
  wire n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2151, n_2152;
  wire n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160;
  wire n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168;
  wire n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178;
  wire n_2179, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187;
  wire n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195;
  wire n_2196, n_2197, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204;
  wire n_2205, n_2206, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214;
  wire n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222;
  wire n_2223, n_2224, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232;
  wire n_2233, n_2234, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241;
  wire n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249;
  wire n_2250, n_2252, n_2253, n_2254, n_2255, n_2257, n_2258, n_2259;
  wire n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268;
  wire n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2277, n_2278;
  wire n_2279, n_2280, n_2281, n_2282, n_2283, n_2285, n_2286, n_2287;
  wire n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295;
  wire n_2296, n_2297, n_2299, n_2301, n_2302, n_2303, n_2304, n_2305;
  wire n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314;
  wire n_2315, n_2316, n_2317, n_2318, n_2321, n_2322, n_2323, n_2324;
  wire n_2325, n_2326, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333;
  wire n_2334, n_2335, n_2336, n_2337, n_2338, n_2340, n_2341, n_2342;
  wire n_2343, n_2345, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352;
  wire n_2353, n_2354, n_2355, n_2356, n_2359, n_2360, n_2361, n_2362;
  wire n_2363, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371;
  wire n_2372, n_2373, n_2375, n_2377, n_2378, n_2379, n_2381, n_2382;
  wire n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2391, n_2392;
  wire n_2393, n_2394, n_2396, n_2397, n_2398, n_2399, n_2400, n_2401;
  wire n_2402, n_2404, n_2406, n_2407, n_2409, n_2410, n_2411, n_2412;
  wire n_2413, n_2414, n_2417, n_2418, n_2419, n_2421, n_2422, n_2423;
  wire n_2424, n_2425, n_2427, n_2428, n_2431, n_2432, n_2433, n_2434;
  wire n_2437, n_2438, n_2440, n_2441, n_2442, n_2445, n_2447, n_2448;
  wire n_2451, n_2453, n_2457, n_2458, n_2459, n_2460, n_2461, n_2462;
  wire n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, n_2469, n_2470;
  wire n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, n_2478;
  wire n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486;
  wire n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, n_2493, n_2494;
  wire n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, n_2502;
  wire n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509, n_2510;
  wire n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517, n_2518;
  wire n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, n_2525, n_2526;
  wire n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, n_2533, n_2534;
  wire n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, n_2542;
  wire n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550;
  wire n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558;
  wire n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, n_2566;
  wire n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574;
  wire n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582;
  wire n_2583, n_2584, n_2585, n_2586, n_2587, n_2588, n_2589, n_2590;
  wire n_2591, n_2592, n_2593, n_2594, n_2595, n_2596, n_2597, n_2598;
  wire n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, n_2606;
  wire n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614;
  wire n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, n_2622;
  wire n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630;
  wire n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, n_2638;
  wire n_2639, n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, n_2646;
  wire n_2647, n_2648, n_2649, n_2650, n_2651, n_2652, n_2653, n_2654;
  wire n_2655, n_2656, n_2657, n_2658, n_2659, n_2660, n_2661, n_2662;
  wire n_2663, n_2664, n_2665, n_2666, n_2667, n_2668, n_2669, n_2670;
  wire n_2671, n_2672, n_2673, n_2674, n_2675, n_2676, n_2677, n_2678;
  wire n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, n_2685, n_2686;
  wire n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2693, n_2694;
  wire n_2695, n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702;
  wire n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, n_2710;
  wire n_2711, n_2712, n_2713, n_2714, n_2715, n_2716, n_2717, n_2718;
  wire n_2719, n_2720, n_2721, n_2722, n_2723, n_2724, n_2725, n_2726;
  wire n_2727, n_2728, n_2729, n_2730, n_2731, n_2732, n_2733, n_2734;
  wire n_2735, n_2736, n_2737, n_2738, n_2739, n_2740, n_2741, n_2742;
  wire n_2743, n_2744, n_2745, n_2746, n_2747, n_2748, n_2749, n_2750;
  wire n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, n_2757, n_2758;
  wire n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, n_2766;
  wire n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774;
  wire n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, n_2781, n_2782;
  wire n_2783, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, n_2790;
  wire n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2798;
  wire n_2799, n_2800, n_2801, n_2802, n_2803, n_2804, n_2805, n_2806;
  wire n_2807, n_2808, n_2809, n_2810, n_2811, n_2812, n_2813, n_2814;
  wire n_2815, n_2816, n_2817, n_2818, n_2819, n_2820, n_2821, n_2822;
  wire n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830;
  wire n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, n_2838;
  wire n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846;
  wire n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, n_2854;
  wire n_2855, n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, n_2862;
  wire n_2863, n_2864, n_2865, n_2866, n_2867, n_2868, n_2869, n_2870;
  wire n_2871, n_2872, n_2873, n_2874, n_2875, n_2876, n_2877, n_2878;
  wire n_2879, n_2880, n_2881, n_2882, n_2883, n_2884, n_2885, n_2886;
  wire n_2887, n_2888, n_2889, n_2890, n_2891, n_2892, n_2893, n_2894;
  wire n_2895, n_2896, n_2897, n_2898, n_2899, n_2900, n_2901, n_2902;
  wire n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2909, n_2910;
  wire n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918;
  wire n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926;
  wire n_2927, n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, n_2934;
  wire n_2935, n_2936, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942;
  wire n_2943, n_2944, n_2945, n_2946, n_2947, n_2948, n_2949, n_2950;
  wire n_2951, n_2952, n_2953, n_2954, n_2955, n_2956, n_2957, n_2958;
  wire n_2959, n_2960, n_2961, n_2962, n_2963, n_2964, n_2965, n_2966;
  wire n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, n_2973, n_2974;
  wire n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, n_2982;
  wire n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990;
  wire n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, n_2997, n_2998;
  wire n_2999, n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, n_3006;
  wire n_3007, n_3008, n_3009, n_3010, n_3011, n_3012, n_3013, n_3014;
  wire n_3015, n_3016, n_3017, n_3018, n_3019, n_3020, n_3021, n_3022;
  wire n_3023, n_3024, n_3025, n_3026, n_3027, n_3028, n_3029, n_3030;
  wire n_3031, n_3032, n_3033, n_3034, n_3035, n_3036, n_3037, n_3038;
  wire n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, n_3045, n_3046;
  wire n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, n_3053, n_3054;
  wire n_3055, n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, n_3062;
  wire n_3063, n_3064, n_3065, n_3066, n_3067, n_3068, n_3069, n_3070;
  wire n_3071, n_3072, n_3073, n_3074, n_3075, n_3076, n_3077, n_3078;
  wire n_3079, n_3080, n_3081, n_3082, n_3083, n_3084, n_3085, n_3086;
  wire n_3087, n_3088, n_3089, n_3090, n_3091, n_3092, n_3093, n_3094;
  wire n_3095, n_3096, n_3097, n_3098, n_3099, n_3100, n_3101, n_3102;
  wire n_3103, n_3104, n_3105, n_3106, n_3107, n_3108, n_3109, n_3110;
  wire n_3111, n_3112, n_3113, n_3114, n_3115, n_3116, n_3117, n_3118;
  wire n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, n_3125, n_3126;
  wire n_3127, n_3128, n_3129, n_3130, n_3131, n_3132, n_3133, n_3134;
  wire n_3135, n_3136, n_3137, n_3138, n_3139, n_3140, n_3141, n_3142;
  wire n_3143, n_3144, n_3145, n_3146, n_3147, n_3148, n_3149, n_3150;
  wire n_3151, n_3152, n_3153, n_3154, n_3155, n_3156, n_3157, n_3158;
  wire n_3159, n_3160, n_3161, n_3162, n_3163, n_3164, n_3165, n_3166;
  wire n_3167, n_3168, n_3169, n_3170, n_3171, n_3172, n_3173, n_3174;
  wire n_3175, n_3176, n_3177, n_3178, n_3179, n_3180, n_3181, n_3182;
  wire n_3183, n_3184, n_3185, n_3186, n_3187, n_3188, n_3189, n_3190;
  wire n_3191, n_3192, n_3193, n_3194, n_3195, n_3196, n_3197, n_3198;
  wire n_3199, n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3206;
  wire n_3207, n_3208, n_3209, n_3210, n_3211, n_3212, n_3213, n_3214;
  wire n_3215, n_3216, n_3217, n_3218, n_3219, n_3220, n_3221, n_3222;
  wire n_3223, n_3224, n_3225, n_3226, n_3227, n_3228, n_3229, n_3230;
  wire n_3231, n_3232, n_3233, n_3234, n_3235, n_3236, n_3237, n_3238;
  wire n_3239, n_3240, n_3241, n_3242, n_3243, n_3244, n_3245, n_3246;
  wire n_3247, n_3248, n_3249, n_3250, n_3251, n_3252, n_3253, n_3254;
  wire n_3255, n_3256, n_3257, n_3258, n_3259, n_3260, n_3261, n_3262;
  wire n_3263, n_3264, n_3265, n_3266, n_3267, n_3268, n_3269, n_3270;
  wire n_3271, n_3272, n_3273, n_3274, n_3275, n_3276, n_3277, n_3278;
  wire n_3279, n_3280, n_3281, n_3282, n_3283, n_3284, n_3285, n_3286;
  wire n_3287, n_3288, n_3289, n_3290, n_3291, n_3292, n_3293, n_3294;
  wire n_3295, n_3296, n_3297, n_3298, n_3299, n_3300, n_3301, n_3302;
  wire n_3303, n_3304, n_3305, n_3306, n_3307, n_3308, n_3309, n_3310;
  wire n_3311, n_3312, n_3313, n_3314, n_3315, n_3316, n_3317, n_3318;
  wire n_3319, n_3320, n_3321, n_3322, n_3323, n_3324, n_3325, n_3326;
  wire n_3327, n_3328, n_3329, n_3330, n_3331, n_3332, n_3333, n_3334;
  wire n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, n_3341, n_3342;
  wire n_3343, n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350;
  wire n_3351, n_3352, n_3353, n_3354, n_3355, n_3356, n_3357, n_3358;
  wire n_3359, n_3360, n_3361, n_3362, n_3363, n_3364, n_3365, n_3366;
  wire n_3367, n_3368, n_3369, n_3370, n_3371, n_3372, n_3373, n_3374;
  wire n_3375, n_3376, n_3377, n_3378, n_3379, n_3380, n_3381, n_3382;
  wire n_3383, n_3384, n_3385, n_3386, n_3387, n_3388, n_3389, n_3390;
  wire n_3391, n_3392, n_3393, n_3394, n_3395, n_3396, n_3397, n_3398;
  wire n_3399, n_3400, n_3401, n_3402, n_3403, n_3404, n_3405, n_3406;
  wire n_3407, n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414;
  wire n_3415, n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422;
  wire n_3423, n_3424, n_3425, n_3426, n_3427, n_3428, n_3429, n_3430;
  wire n_3431, n_3432, n_3433, n_3434, n_3435, n_3436, n_3437, n_3438;
  wire n_3439, n_3440, n_3441, n_3442, n_3443, n_3444, n_3445, n_3446;
  wire n_3447, n_3448, n_3449, n_3450, n_3451, n_3452, n_3453, n_3454;
  wire n_3455, n_3456, n_3457, n_3458, n_3459, n_3460, n_3461, n_3462;
  wire n_3463, n_3464, n_3465, n_3466, n_3467, n_3468, n_3469, n_3470;
  wire n_3471, n_3472, n_3473, n_3474, n_3475, n_3476, n_3477, n_3478;
  wire n_3479, n_3480, n_3481, n_3482, n_3483, n_3484, n_3485, n_3486;
  wire n_3487, n_3488, n_3489, n_3490, n_3491, n_3492, n_3493, n_3494;
  wire n_3495, n_3496, n_3497, n_3498, n_3499, n_3500, n_3501, n_3502;
  wire n_3503, n_3504, n_3505, n_3506, n_3507, n_3508, n_3530, n_3533;
  wire n_3535, n_3536, n_3537, n_3538, n_3539, n_3541, n_3542, n_3543;
  wire n_3544, n_3545, n_3547, n_3548, n_3549, n_3550, n_3551, n_3553;
  wire n_3554, n_3555, n_3556, n_3557, n_3559, n_3560, n_3561, n_3562;
  wire n_3563, n_3565, n_3566, n_3567, n_3568, n_3569, n_3571, n_3572;
  wire n_3573, n_3574, n_3575, n_3577, n_3578, n_3579, n_3580, n_3581;
  wire n_3583, n_3584, n_3585, n_3586, n_3587, n_3589, n_3590, n_3591;
  wire n_3592, n_3593, n_3595, n_3596, n_3597, n_3598, n_3599, n_3601;
  wire n_3602, n_3603, n_3604, n_3605, n_3607, n_3608, n_3609, n_3610;
  wire n_3611, n_3613, n_3614, n_3615, n_3616, n_3617, n_3619, n_3620;
  wire n_3621, n_3622, n_3623, n_3625, n_3626, n_3627, n_3628, n_3629;
  wire n_3631, n_3632, n_3633, n_3634, n_3635, n_3637, n_3638, n_3639;
  wire n_3640, n_3641, n_3643, n_3644, n_3645, n_3646, n_3647, n_3649;
  wire n_3650, n_3651, n_3652, n_3653, n_3655, n_3656, n_3657, n_3658;
  wire n_3659, n_3661, n_3662, n_3663, n_3664, n_3665, n_3667, n_3668;
  wire n_3669, n_3670, n_3671, n_3679, n_3683, n_3685, n_3686, n_3688;
  wire n_3689, n_3691, n_3693, n_3695, n_3696, n_3698, n_3699, n_3701;
  wire n_3703, n_3705, n_3706, n_3708, n_3709, n_3711, n_3713, n_3715;
  wire n_3716, n_3718, n_3719, n_3721, n_3723, n_3725, n_3726, n_3728;
  wire n_3729, n_3731, n_3733, n_3735, n_3736, n_3738, n_3739, n_3741;
  wire n_3743, n_3745, n_3746, n_3748, n_3749, n_3751, n_3753, n_3755;
  wire n_3756, n_3758, n_3759, n_3761, n_3763, n_3765, n_3766, n_3768;
  wire n_3769, n_3771, n_3773, n_3775, n_3776, n_3778, n_3779, n_3781;
  wire n_3783, n_3785, n_3786, n_3788, n_3789, n_3791, n_3799, n_3803;
  wire n_3805, n_3806, n_3808, n_3810, n_3812, n_3813, n_3814, n_3816;
  wire n_3817, n_3818, n_3820, n_3821, n_3823, n_3825, n_3827, n_3828;
  wire n_3829, n_3831, n_3832, n_3833, n_3835, n_3836, n_3838, n_3840;
  wire n_3842, n_3843, n_3844, n_3846, n_3847, n_3848, n_3850, n_3851;
  wire n_3853, n_3855, n_3857, n_3858, n_3859, n_3861, n_3862, n_3863;
  wire n_3865, n_3866, n_3868, n_3870, n_3872, n_3873, n_3874, n_3876;
  wire n_3877, n_3878, n_3882, n_3883, n_3884, n_3886, n_3887, n_3889;
  wire n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3896, n_3897;
  wire n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, n_3905, n_3908;
  wire n_3910, n_3911, n_3912, n_3915, n_3918, n_3920, n_3921, n_3923;
  wire n_3925, n_3926, n_3928, n_3930, n_3931, n_3933, n_3935, n_3936;
  wire n_3938, n_3939, n_3941, n_3944, n_3946, n_3947, n_3948, n_3951;
  wire n_3954, n_3956, n_3957, n_3959, n_3961, n_3962, n_3964, n_3966;
  wire n_3967, n_3969, n_3971, n_3972, n_3974, n_3976, n_3977, n_3978;
  wire n_3980, n_3981, n_3983, n_3984, n_3985, n_3986, n_3987, n_3988;
  wire n_3989, n_3990, n_3991, n_3992, n_3993, n_3994, n_3996, n_3997;
  wire n_3998, n_4000, n_4001, n_4002, n_4004, n_4005, n_4006, n_4008;
  wire n_4009, n_4010, n_4012, n_4013, n_4014, n_4016, n_4017, n_4018;
  wire n_4020, n_4021, n_4022, n_4024, n_4025, n_4026, n_4027, n_4029;
  wire n_4031, n_4033, n_4034, n_4035, n_4037, n_4039, n_4040, n_4041;
  wire n_4043, n_4044, n_4046, n_4047, n_4048, n_4049, n_4050, n_4051;
  wire n_4052, n_4053, n_4054, n_4055, n_4056, n_4057, n_4059, n_4060;
  wire n_4061, n_4063, n_4064, n_4065, n_4067, n_4068, n_4069, n_4071;
  wire n_4072, n_4073, n_4075, n_4076, n_4077, n_4079, n_4080, n_4081;
  wire n_4083, n_4084, n_4086, n_4087, n_4088, n_4089, n_4090, n_4091;
  wire n_4092, n_4093, n_4094, n_4095, n_4101, n_4106, n_4109, n_4110;
  wire n_4112, n_4113, n_4114, n_4115, n_4117, n_4118, n_4120, n_4121;
  wire n_4123, n_4124, n_4125, n_4126, n_4128, n_4129, n_4130, n_4132;
  wire n_4133, n_4134, n_4135, n_4137, n_4138, n_4140, n_4141, n_4143;
  wire n_4144, n_4145, n_4146, n_4148, n_4149, n_4150, n_4151, n_4153;
  wire n_4154, n_4155, n_4156, n_4158, n_4159, n_4161, n_4162, n_4164;
  wire n_4165, n_4166, n_4167, n_4169, n_4170, n_4171, n_4173, n_4174;
  wire n_4175, n_4176, n_4178, n_4179, n_4181, n_4182, n_4184, n_4185;
  wire n_4186, n_4187, n_4189, n_4190, n_4191, n_4192, n_4194, n_4195;
  wire n_4196, n_4197, n_4199, n_4200, n_4202, n_4203, n_4205, n_4206;
  wire n_4207, n_4208, n_4210, n_4211, n_4213, n_4214, n_4216, n_4217;
  wire n_4218, n_4219, n_4221, n_4222;
  assign Z[0] = 1'b0;
  assign Z[1] = 1'b0;
  assign Z[2] = 1'b0;
  assign Z[3] = 1'b0;
  xor g126 (n_311, B[2], B[1]);
  xor g127 (n_313, B[3], B[2]);
  nor g131 (n_406, B[1], B[2]);
  nand g132 (n_404, B[1], B[2]);
  xor g138 (n_319, B[3], A[1]);
  xor g142 (n_322, B[3], A[2]);
  nand g143 (n_323, n_322, n_311);
  nand g144 (n_324, n_319, n_315);
  nand g145 (n_204, n_323, n_324);
  xor g146 (n_325, B[3], A[3]);
  nand g147 (n_326, n_325, n_311);
  nand g148 (n_327, n_322, n_315);
  nand g149 (n_151, n_326, n_327);
  xor g150 (n_328, B[3], A[4]);
  nand g151 (n_329, n_328, n_311);
  nand g152 (n_330, n_325, n_315);
  nand g153 (n_150, n_329, n_330);
  xor g154 (n_331, B[3], A[5]);
  nand g155 (n_332, n_331, n_311);
  nand g156 (n_333, n_328, n_315);
  nand g157 (n_1599, n_332, n_333);
  xor g158 (n_334, B[3], A[6]);
  nand g159 (n_335, n_334, n_311);
  nand g160 (n_336, n_331, n_315);
  nand g161 (n_1603, n_335, n_336);
  xor g162 (n_337, B[3], A[7]);
  nand g163 (n_338, n_337, n_311);
  nand g164 (n_339, n_334, n_315);
  nand g165 (n_1607, n_338, n_339);
  xor g166 (n_340, B[3], A[8]);
  nand g167 (n_341, n_340, n_311);
  nand g168 (n_342, n_337, n_315);
  nand g169 (n_1613, n_341, n_342);
  xor g170 (n_343, B[3], A[9]);
  nand g171 (n_344, n_343, n_311);
  nand g172 (n_345, n_340, n_315);
  nand g173 (n_1622, n_344, n_345);
  xor g174 (n_346, B[3], A[10]);
  nand g175 (n_347, n_346, n_311);
  nand g176 (n_348, n_343, n_315);
  nand g177 (n_1632, n_347, n_348);
  xor g178 (n_349, B[3], A[11]);
  nand g179 (n_350, n_349, n_311);
  nand g180 (n_351, n_346, n_315);
  nand g181 (n_1641, n_350, n_351);
  xor g182 (n_352, B[3], A[12]);
  nand g183 (n_353, n_352, n_311);
  nand g184 (n_354, n_349, n_315);
  nand g185 (n_1655, n_353, n_354);
  xor g186 (n_355, B[3], A[13]);
  nand g187 (n_356, n_355, n_311);
  nand g188 (n_357, n_352, n_315);
  nand g189 (n_1668, n_356, n_357);
  xor g190 (n_358, B[3], A[14]);
  nand g191 (n_359, n_358, n_311);
  nand g192 (n_360, n_355, n_315);
  nand g193 (n_1684, n_359, n_360);
  xor g194 (n_361, B[3], A[15]);
  nand g195 (n_362, n_361, n_311);
  nand g196 (n_363, n_358, n_315);
  nand g197 (n_1700, n_362, n_363);
  xor g198 (n_364, B[3], A[16]);
  nand g199 (n_365, n_364, n_311);
  nand g200 (n_366, n_361, n_315);
  nand g201 (n_1715, n_365, n_366);
  xor g202 (n_367, B[3], A[17]);
  nand g203 (n_368, n_367, n_311);
  nand g204 (n_369, n_364, n_315);
  nand g205 (n_1732, n_368, n_369);
  xor g206 (n_370, B[3], A[18]);
  nand g207 (n_371, n_370, n_311);
  nand g208 (n_372, n_367, n_315);
  nand g209 (n_1754, n_371, n_372);
  xor g210 (n_373, B[3], A[19]);
  nand g211 (n_374, n_373, n_311);
  nand g212 (n_375, n_370, n_315);
  nand g213 (n_1777, n_374, n_375);
  xor g214 (n_376, B[3], A[20]);
  nand g215 (n_377, n_376, n_311);
  nand g216 (n_378, n_373, n_315);
  nand g217 (n_1798, n_377, n_378);
  xor g218 (n_379, B[3], A[21]);
  nand g219 (n_380, n_379, n_311);
  nand g220 (n_381, n_376, n_315);
  nand g221 (n_1827, n_380, n_381);
  xor g222 (n_382, B[3], A[22]);
  nand g223 (n_383, n_382, n_311);
  nand g224 (n_384, n_379, n_315);
  nand g225 (n_1850, n_383, n_384);
  xor g226 (n_385, B[3], A[23]);
  nand g227 (n_386, n_385, n_311);
  nand g228 (n_387, n_382, n_315);
  nand g229 (n_1882, n_386, n_387);
  xor g230 (n_388, B[3], A[24]);
  nand g231 (n_389, n_388, n_311);
  nand g232 (n_390, n_385, n_315);
  nand g233 (n_1914, n_389, n_390);
  xor g234 (n_391, B[3], A[25]);
  nand g235 (n_392, n_391, n_311);
  nand g236 (n_393, n_388, n_315);
  nand g237 (n_1949, n_392, n_393);
  nand g239 (n_396, B[3], n_311);
  nand g240 (n_397, n_391, n_315);
  nand g241 (n_1973, n_396, n_397);
  nand g244 (n_401, B[3], n_315);
  nand g245 (n_402, n_396, n_401);
  or g249 (n_407, n_405, n_406);
  and g250 (n_152, B[3], n_407);
  xor g251 (n_408, B[4], B[3]);
  xor g252 (n_410, B[5], B[4]);
  nor g256 (n_503, B[3], B[4]);
  nand g257 (n_501, B[3], B[4]);
  xor g263 (n_416, B[5], A[1]);
  xor g267 (n_419, B[5], A[2]);
  nand g268 (n_420, n_419, n_408);
  nand g269 (n_421, n_416, n_412);
  nand g270 (n_1598, n_420, n_421);
  xor g271 (n_422, B[5], A[3]);
  nand g272 (n_423, n_422, n_408);
  nand g273 (n_424, n_419, n_412);
  nand g274 (n_1600, n_423, n_424);
  xor g275 (n_425, B[5], A[4]);
  nand g276 (n_426, n_425, n_408);
  nand g277 (n_427, n_422, n_412);
  nand g278 (n_1602, n_426, n_427);
  xor g279 (n_428, B[5], A[5]);
  nand g280 (n_429, n_428, n_408);
  nand g281 (n_430, n_425, n_412);
  nand g282 (n_1608, n_429, n_430);
  xor g283 (n_431, B[5], A[6]);
  nand g284 (n_432, n_431, n_408);
  nand g285 (n_433, n_428, n_412);
  nand g286 (n_1612, n_432, n_433);
  xor g287 (n_434, B[5], A[7]);
  nand g288 (n_435, n_434, n_408);
  nand g289 (n_436, n_431, n_412);
  nand g290 (n_1621, n_435, n_436);
  xor g291 (n_437, B[5], A[8]);
  nand g292 (n_438, n_437, n_408);
  nand g293 (n_439, n_434, n_412);
  nand g294 (n_1628, n_438, n_439);
  xor g295 (n_440, B[5], A[9]);
  nand g296 (n_441, n_440, n_408);
  nand g297 (n_442, n_437, n_412);
  nand g298 (n_1640, n_441, n_442);
  xor g299 (n_443, B[5], A[10]);
  nand g300 (n_444, n_443, n_408);
  nand g301 (n_445, n_440, n_412);
  nand g302 (n_1650, n_444, n_445);
  xor g303 (n_446, B[5], A[11]);
  nand g304 (n_447, n_446, n_408);
  nand g305 (n_448, n_443, n_412);
  nand g306 (n_1664, n_447, n_448);
  xor g307 (n_449, B[5], A[12]);
  nand g308 (n_450, n_449, n_408);
  nand g309 (n_451, n_446, n_412);
  nand g310 (n_1679, n_450, n_451);
  xor g311 (n_452, B[5], A[13]);
  nand g312 (n_453, n_452, n_408);
  nand g313 (n_454, n_449, n_412);
  nand g314 (n_1698, n_453, n_454);
  xor g315 (n_455, B[5], A[14]);
  nand g316 (n_456, n_455, n_408);
  nand g317 (n_457, n_452, n_412);
  nand g318 (n_1719, n_456, n_457);
  xor g319 (n_458, B[5], A[15]);
  nand g320 (n_459, n_458, n_408);
  nand g321 (n_460, n_455, n_412);
  nand g322 (n_1735, n_459, n_460);
  xor g323 (n_461, B[5], A[16]);
  nand g324 (n_462, n_461, n_408);
  nand g325 (n_463, n_458, n_412);
  nand g326 (n_1757, n_462, n_463);
  xor g327 (n_464, B[5], A[17]);
  nand g328 (n_465, n_464, n_408);
  nand g329 (n_466, n_461, n_412);
  nand g330 (n_1775, n_465, n_466);
  xor g331 (n_467, B[5], A[18]);
  nand g332 (n_468, n_467, n_408);
  nand g333 (n_469, n_464, n_412);
  nand g334 (n_1800, n_468, n_469);
  xor g335 (n_470, B[5], A[19]);
  nand g336 (n_471, n_470, n_408);
  nand g337 (n_472, n_467, n_412);
  nand g338 (n_1830, n_471, n_472);
  xor g339 (n_473, B[5], A[20]);
  nand g340 (n_474, n_473, n_408);
  nand g341 (n_475, n_470, n_412);
  nand g342 (n_1858, n_474, n_475);
  xor g343 (n_476, B[5], A[21]);
  nand g344 (n_477, n_476, n_408);
  nand g345 (n_478, n_473, n_412);
  nand g346 (n_1886, n_477, n_478);
  xor g347 (n_479, B[5], A[22]);
  nand g348 (n_480, n_479, n_408);
  nand g349 (n_481, n_476, n_412);
  nand g350 (n_1916, n_480, n_481);
  xor g351 (n_482, B[5], A[23]);
  nand g352 (n_483, n_482, n_408);
  nand g353 (n_484, n_479, n_412);
  nand g354 (n_1948, n_483, n_484);
  xor g355 (n_485, B[5], A[24]);
  nand g356 (n_486, n_485, n_408);
  nand g357 (n_487, n_482, n_412);
  nand g358 (n_1982, n_486, n_487);
  xor g359 (n_488, B[5], A[25]);
  nand g360 (n_489, n_488, n_408);
  nand g361 (n_490, n_485, n_412);
  nand g362 (n_2013, n_489, n_490);
  nand g364 (n_493, B[5], n_408);
  nand g365 (n_494, n_488, n_412);
  nand g366 (n_2042, n_493, n_494);
  nand g369 (n_498, B[5], n_412);
  nand g370 (n_499, n_493, n_498);
  or g374 (n_504, n_502, n_503);
  and g375 (n_1597, B[5], n_504);
  xor g376 (n_505, B[6], B[5]);
  xor g377 (n_507, B[7], B[6]);
  nor g381 (n_600, B[5], B[6]);
  nand g382 (n_598, B[5], B[6]);
  xor g388 (n_513, B[7], A[1]);
  xor g392 (n_516, B[7], A[2]);
  nand g393 (n_517, n_516, n_505);
  nand g394 (n_518, n_513, n_509);
  nand g395 (n_1604, n_517, n_518);
  xor g396 (n_519, B[7], A[3]);
  nand g397 (n_520, n_519, n_505);
  nand g398 (n_521, n_516, n_509);
  nand g399 (n_1606, n_520, n_521);
  xor g400 (n_522, B[7], A[4]);
  nand g401 (n_523, n_522, n_505);
  nand g402 (n_524, n_519, n_509);
  nand g403 (n_1615, n_523, n_524);
  xor g404 (n_525, B[7], A[5]);
  nand g405 (n_526, n_525, n_505);
  nand g406 (n_527, n_522, n_509);
  nand g407 (n_1620, n_526, n_527);
  xor g408 (n_528, B[7], A[6]);
  nand g409 (n_529, n_528, n_505);
  nand g410 (n_530, n_525, n_509);
  nand g411 (n_1630, n_529, n_530);
  xor g412 (n_531, B[7], A[7]);
  nand g413 (n_532, n_531, n_505);
  nand g414 (n_533, n_528, n_509);
  nand g415 (n_1639, n_532, n_533);
  xor g416 (n_534, B[7], A[8]);
  nand g417 (n_535, n_534, n_505);
  nand g418 (n_536, n_531, n_509);
  nand g419 (n_1653, n_535, n_536);
  xor g420 (n_537, B[7], A[9]);
  nand g421 (n_538, n_537, n_505);
  nand g422 (n_539, n_534, n_509);
  nand g423 (n_1667, n_538, n_539);
  xor g424 (n_540, B[7], A[10]);
  nand g425 (n_541, n_540, n_505);
  nand g426 (n_542, n_537, n_509);
  nand g427 (n_1683, n_541, n_542);
  xor g428 (n_543, B[7], A[11]);
  nand g429 (n_544, n_543, n_505);
  nand g430 (n_545, n_540, n_509);
  nand g431 (n_1695, n_544, n_545);
  xor g432 (n_546, B[7], A[12]);
  nand g433 (n_547, n_546, n_505);
  nand g434 (n_548, n_543, n_509);
  nand g435 (n_1713, n_547, n_548);
  xor g436 (n_549, B[7], A[13]);
  nand g437 (n_550, n_549, n_505);
  nand g438 (n_551, n_546, n_509);
  nand g439 (n_1736, n_550, n_551);
  xor g440 (n_552, B[7], A[14]);
  nand g441 (n_553, n_552, n_505);
  nand g442 (n_554, n_549, n_509);
  nand g443 (n_1758, n_553, n_554);
  xor g444 (n_555, B[7], A[15]);
  nand g445 (n_556, n_555, n_505);
  nand g446 (n_557, n_552, n_509);
  nand g447 (n_1779, n_556, n_557);
  xor g448 (n_558, B[7], A[16]);
  nand g449 (n_559, n_558, n_505);
  nand g450 (n_560, n_555, n_509);
  nand g451 (n_1803, n_559, n_560);
  xor g452 (n_561, B[7], A[17]);
  nand g453 (n_562, n_561, n_505);
  nand g454 (n_563, n_558, n_509);
  nand g455 (n_1831, n_562, n_563);
  xor g456 (n_564, B[7], A[18]);
  nand g457 (n_565, n_564, n_505);
  nand g458 (n_566, n_561, n_509);
  nand g459 (n_1859, n_565, n_566);
  xor g460 (n_567, B[7], A[19]);
  nand g461 (n_568, n_567, n_505);
  nand g462 (n_569, n_564, n_509);
  nand g463 (n_1881, n_568, n_569);
  xor g464 (n_570, B[7], A[20]);
  nand g465 (n_571, n_570, n_505);
  nand g466 (n_572, n_567, n_509);
  nand g467 (n_1912, n_571, n_572);
  xor g468 (n_573, B[7], A[21]);
  nand g469 (n_574, n_573, n_505);
  nand g470 (n_575, n_570, n_509);
  nand g471 (n_1944, n_574, n_575);
  xor g472 (n_576, B[7], A[22]);
  nand g473 (n_577, n_576, n_505);
  nand g474 (n_578, n_573, n_509);
  nand g475 (n_1980, n_577, n_578);
  xor g476 (n_579, B[7], A[23]);
  nand g477 (n_580, n_579, n_505);
  nand g478 (n_581, n_576, n_509);
  nand g479 (n_2010, n_580, n_581);
  xor g480 (n_582, B[7], A[24]);
  nand g481 (n_583, n_582, n_505);
  nand g482 (n_584, n_579, n_509);
  nand g483 (n_2047, n_583, n_584);
  xor g484 (n_585, B[7], A[25]);
  nand g485 (n_586, n_585, n_505);
  nand g486 (n_587, n_582, n_509);
  nand g487 (n_2081, n_586, n_587);
  nand g489 (n_590, B[7], n_505);
  nand g490 (n_591, n_585, n_509);
  nand g491 (n_2114, n_590, n_591);
  nand g494 (n_595, B[7], n_509);
  nand g495 (n_596, n_590, n_595);
  or g499 (n_601, n_599, n_600);
  and g500 (n_1601, B[7], n_601);
  xor g501 (n_602, B[8], B[7]);
  xor g502 (n_604, B[9], B[8]);
  nor g506 (n_697, B[7], B[8]);
  nand g507 (n_695, B[7], B[8]);
  xor g513 (n_610, B[9], A[1]);
  xor g517 (n_613, B[9], A[2]);
  nand g518 (n_614, n_613, n_602);
  nand g519 (n_615, n_610, n_606);
  nand g520 (n_1614, n_614, n_615);
  xor g521 (n_616, B[9], A[3]);
  nand g522 (n_617, n_616, n_602);
  nand g523 (n_618, n_613, n_606);
  nand g524 (n_1619, n_617, n_618);
  xor g525 (n_619, B[9], A[4]);
  nand g526 (n_620, n_619, n_602);
  nand g527 (n_621, n_616, n_606);
  nand g528 (n_1629, n_620, n_621);
  xor g529 (n_622, B[9], A[5]);
  nand g530 (n_623, n_622, n_602);
  nand g531 (n_624, n_619, n_606);
  nand g532 (n_1642, n_623, n_624);
  xor g533 (n_625, B[9], A[6]);
  nand g534 (n_626, n_625, n_602);
  nand g535 (n_627, n_622, n_606);
  nand g536 (n_1654, n_626, n_627);
  xor g537 (n_628, B[9], A[7]);
  nand g538 (n_629, n_628, n_602);
  nand g539 (n_630, n_625, n_606);
  nand g540 (n_1666, n_629, n_630);
  xor g541 (n_631, B[9], A[8]);
  nand g542 (n_632, n_631, n_602);
  nand g543 (n_633, n_628, n_606);
  nand g544 (n_1678, n_632, n_633);
  xor g545 (n_634, B[9], A[9]);
  nand g546 (n_635, n_634, n_602);
  nand g547 (n_636, n_631, n_606);
  nand g548 (n_1697, n_635, n_636);
  xor g549 (n_637, B[9], A[10]);
  nand g550 (n_638, n_637, n_602);
  nand g551 (n_639, n_634, n_606);
  nand g552 (n_1716, n_638, n_639);
  xor g553 (n_640, B[9], A[11]);
  nand g554 (n_641, n_640, n_602);
  nand g555 (n_642, n_637, n_606);
  nand g556 (n_1737, n_641, n_642);
  xor g557 (n_643, B[9], A[12]);
  nand g558 (n_644, n_643, n_602);
  nand g559 (n_645, n_640, n_606);
  nand g560 (n_1759, n_644, n_645);
  xor g561 (n_646, B[9], A[13]);
  nand g562 (n_647, n_646, n_602);
  nand g563 (n_648, n_643, n_606);
  nand g564 (n_1780, n_647, n_648);
  xor g565 (n_649, B[9], A[14]);
  nand g566 (n_650, n_649, n_602);
  nand g567 (n_651, n_646, n_606);
  nand g568 (n_1805, n_650, n_651);
  xor g569 (n_652, B[9], A[15]);
  nand g570 (n_653, n_652, n_602);
  nand g571 (n_654, n_649, n_606);
  nand g572 (n_1828, n_653, n_654);
  xor g573 (n_655, B[9], A[16]);
  nand g574 (n_656, n_655, n_602);
  nand g575 (n_657, n_652, n_606);
  nand g576 (n_1856, n_656, n_657);
  xor g577 (n_658, B[9], A[17]);
  nand g578 (n_659, n_658, n_602);
  nand g579 (n_660, n_655, n_606);
  nand g580 (n_1887, n_659, n_660);
  xor g581 (n_661, B[9], A[18]);
  nand g582 (n_662, n_661, n_602);
  nand g583 (n_663, n_658, n_606);
  nand g584 (n_1917, n_662, n_663);
  xor g585 (n_664, B[9], A[19]);
  nand g586 (n_665, n_664, n_602);
  nand g587 (n_666, n_661, n_606);
  nand g588 (n_1943, n_665, n_666);
  xor g589 (n_667, B[9], A[20]);
  nand g590 (n_668, n_667, n_602);
  nand g591 (n_669, n_664, n_606);
  nand g592 (n_1977, n_668, n_669);
  xor g593 (n_670, B[9], A[21]);
  nand g594 (n_671, n_670, n_602);
  nand g595 (n_672, n_667, n_606);
  nand g596 (n_2008, n_671, n_672);
  xor g597 (n_673, B[9], A[22]);
  nand g598 (n_674, n_673, n_602);
  nand g599 (n_675, n_670, n_606);
  nand g600 (n_2046, n_674, n_675);
  xor g601 (n_676, B[9], A[23]);
  nand g602 (n_677, n_676, n_602);
  nand g603 (n_678, n_673, n_606);
  nand g604 (n_2076, n_677, n_678);
  xor g605 (n_679, B[9], A[24]);
  nand g606 (n_680, n_679, n_602);
  nand g607 (n_681, n_676, n_606);
  nand g608 (n_2110, n_680, n_681);
  xor g609 (n_682, B[9], A[25]);
  nand g610 (n_683, n_682, n_602);
  nand g611 (n_684, n_679, n_606);
  nand g612 (n_2141, n_683, n_684);
  nand g614 (n_687, B[9], n_602);
  nand g615 (n_688, n_682, n_606);
  nand g616 (n_2177, n_687, n_688);
  nand g619 (n_692, B[9], n_606);
  nand g620 (n_693, n_687, n_692);
  or g624 (n_698, n_696, n_697);
  and g625 (n_1611, B[9], n_698);
  xor g626 (n_699, B[10], B[9]);
  xor g627 (n_701, B[11], B[10]);
  nor g631 (n_794, B[9], B[10]);
  nand g632 (n_792, B[9], B[10]);
  xor g638 (n_707, B[11], A[1]);
  xor g642 (n_710, B[11], A[2]);
  nand g643 (n_711, n_710, n_699);
  nand g644 (n_712, n_707, n_703);
  nand g645 (n_1631, n_711, n_712);
  xor g646 (n_713, B[11], A[3]);
  nand g647 (n_714, n_713, n_699);
  nand g648 (n_715, n_710, n_703);
  nand g649 (n_1638, n_714, n_715);
  xor g650 (n_716, B[11], A[4]);
  nand g651 (n_717, n_716, n_699);
  nand g652 (n_718, n_713, n_703);
  nand g653 (n_1651, n_717, n_718);
  xor g654 (n_719, B[11], A[5]);
  nand g655 (n_720, n_719, n_699);
  nand g656 (n_721, n_716, n_703);
  nand g657 (n_1665, n_720, n_721);
  xor g658 (n_722, B[11], A[6]);
  nand g659 (n_723, n_722, n_699);
  nand g660 (n_724, n_719, n_703);
  nand g661 (n_1680, n_723, n_724);
  xor g662 (n_725, B[11], A[7]);
  nand g663 (n_726, n_725, n_699);
  nand g664 (n_727, n_722, n_703);
  nand g665 (n_1699, n_726, n_727);
  xor g666 (n_728, B[11], A[8]);
  nand g667 (n_729, n_728, n_699);
  nand g668 (n_730, n_725, n_703);
  nand g669 (n_1712, n_729, n_730);
  xor g670 (n_731, B[11], A[9]);
  nand g671 (n_732, n_731, n_699);
  nand g672 (n_733, n_728, n_703);
  nand g673 (n_1734, n_732, n_733);
  xor g674 (n_734, B[11], A[10]);
  nand g675 (n_735, n_734, n_699);
  nand g676 (n_736, n_731, n_703);
  nand g677 (n_1756, n_735, n_736);
  xor g678 (n_737, B[11], A[11]);
  nand g679 (n_738, n_737, n_699);
  nand g680 (n_739, n_734, n_703);
  nand g681 (n_1781, n_738, n_739);
  xor g682 (n_740, B[11], A[12]);
  nand g683 (n_741, n_740, n_699);
  nand g684 (n_742, n_737, n_703);
  nand g685 (n_1806, n_741, n_742);
  xor g686 (n_743, B[11], A[13]);
  nand g687 (n_744, n_743, n_699);
  nand g688 (n_745, n_740, n_703);
  nand g689 (n_1826, n_744, n_745);
  xor g690 (n_746, B[11], A[14]);
  nand g691 (n_747, n_746, n_699);
  nand g692 (n_748, n_743, n_703);
  nand g693 (n_1854, n_747, n_748);
  xor g694 (n_749, B[11], A[15]);
  nand g695 (n_750, n_749, n_699);
  nand g696 (n_751, n_746, n_703);
  nand g697 (n_1883, n_750, n_751);
  xor g698 (n_752, B[11], A[16]);
  nand g699 (n_753, n_752, n_699);
  nand g700 (n_754, n_749, n_703);
  nand g701 (n_1915, n_753, n_754);
  xor g702 (n_755, B[11], A[17]);
  nand g703 (n_756, n_755, n_699);
  nand g704 (n_757, n_752, n_703);
  nand g705 (n_1942, n_756, n_757);
  xor g706 (n_758, B[11], A[18]);
  nand g707 (n_759, n_758, n_699);
  nand g708 (n_760, n_755, n_703);
  nand g709 (n_1983, n_759, n_760);
  xor g710 (n_761, B[11], A[19]);
  nand g711 (n_762, n_761, n_699);
  nand g712 (n_763, n_758, n_703);
  nand g713 (n_2017, n_762, n_763);
  xor g714 (n_764, B[11], A[20]);
  nand g715 (n_765, n_764, n_699);
  nand g716 (n_766, n_761, n_703);
  nand g717 (n_2051, n_765, n_766);
  xor g718 (n_767, B[11], A[21]);
  nand g719 (n_768, n_767, n_699);
  nand g720 (n_769, n_764, n_703);
  nand g721 (n_2085, n_768, n_769);
  xor g722 (n_770, B[11], A[22]);
  nand g723 (n_771, n_770, n_699);
  nand g724 (n_772, n_767, n_703);
  nand g725 (n_2116, n_771, n_772);
  xor g726 (n_773, B[11], A[23]);
  nand g727 (n_774, n_773, n_699);
  nand g728 (n_775, n_770, n_703);
  nand g729 (n_2149, n_774, n_775);
  xor g730 (n_776, B[11], A[24]);
  nand g731 (n_777, n_776, n_699);
  nand g732 (n_778, n_773, n_703);
  nand g733 (n_2179, n_777, n_778);
  xor g734 (n_779, B[11], A[25]);
  nand g735 (n_780, n_779, n_699);
  nand g736 (n_781, n_776, n_703);
  nand g737 (n_2204, n_780, n_781);
  nand g739 (n_784, B[11], n_699);
  nand g740 (n_785, n_779, n_703);
  nand g741 (n_2227, n_784, n_785);
  nand g744 (n_789, B[11], n_703);
  nand g745 (n_790, n_784, n_789);
  or g749 (n_795, n_793, n_794);
  and g750 (n_1627, B[11], n_795);
  xor g751 (n_796, B[12], B[11]);
  xor g752 (n_798, B[13], B[12]);
  nor g756 (n_891, B[11], B[12]);
  nand g757 (n_889, B[11], B[12]);
  xor g763 (n_804, B[13], A[1]);
  xor g767 (n_807, B[13], A[2]);
  nand g768 (n_808, n_807, n_796);
  nand g769 (n_809, n_804, n_800);
  nand g770 (n_1652, n_808, n_809);
  xor g771 (n_810, B[13], A[3]);
  nand g772 (n_811, n_810, n_796);
  nand g773 (n_812, n_807, n_800);
  nand g774 (n_1663, n_811, n_812);
  xor g775 (n_813, B[13], A[4]);
  nand g776 (n_814, n_813, n_796);
  nand g777 (n_815, n_810, n_800);
  nand g778 (n_1682, n_814, n_815);
  xor g779 (n_816, B[13], A[5]);
  nand g780 (n_817, n_816, n_796);
  nand g781 (n_818, n_813, n_800);
  nand g782 (n_1696, n_817, n_818);
  xor g783 (n_819, B[13], A[6]);
  nand g784 (n_820, n_819, n_796);
  nand g785 (n_821, n_816, n_800);
  nand g786 (n_1714, n_820, n_821);
  xor g787 (n_822, B[13], A[7]);
  nand g788 (n_823, n_822, n_796);
  nand g789 (n_824, n_819, n_800);
  nand g790 (n_1738, n_823, n_824);
  xor g791 (n_825, B[13], A[8]);
  nand g792 (n_826, n_825, n_796);
  nand g793 (n_827, n_822, n_800);
  nand g794 (n_1752, n_826, n_827);
  xor g795 (n_828, B[13], A[9]);
  nand g796 (n_829, n_828, n_796);
  nand g797 (n_830, n_825, n_800);
  nand g798 (n_1778, n_829, n_830);
  xor g799 (n_831, B[13], A[10]);
  nand g800 (n_832, n_831, n_796);
  nand g801 (n_833, n_828, n_800);
  nand g802 (n_1804, n_832, n_833);
  xor g803 (n_834, B[13], A[11]);
  nand g804 (n_835, n_834, n_796);
  nand g805 (n_836, n_831, n_800);
  nand g806 (n_1824, n_835, n_836);
  xor g807 (n_837, B[13], A[12]);
  nand g808 (n_838, n_837, n_796);
  nand g809 (n_839, n_834, n_800);
  nand g810 (n_1855, n_838, n_839);
  xor g811 (n_840, B[13], A[13]);
  nand g812 (n_841, n_840, n_796);
  nand g813 (n_842, n_837, n_800);
  nand g814 (n_1884, n_841, n_842);
  xor g815 (n_843, B[13], A[14]);
  nand g816 (n_844, n_843, n_796);
  nand g817 (n_845, n_840, n_800);
  nand g818 (n_1908, n_844, n_845);
  xor g819 (n_846, B[13], A[15]);
  nand g820 (n_847, n_846, n_796);
  nand g821 (n_848, n_843, n_800);
  nand g822 (n_1945, n_847, n_848);
  xor g823 (n_849, B[13], A[16]);
  nand g824 (n_850, n_849, n_796);
  nand g825 (n_851, n_846, n_800);
  nand g826 (n_1974, n_850, n_851);
  xor g827 (n_852, B[13], A[17]);
  nand g828 (n_853, n_852, n_796);
  nand g829 (n_854, n_849, n_800);
  nand g830 (n_2006, n_853, n_854);
  xor g831 (n_855, B[13], A[18]);
  nand g832 (n_856, n_855, n_796);
  nand g833 (n_857, n_852, n_800);
  nand g834 (n_2050, n_856, n_857);
  xor g835 (n_858, B[13], A[19]);
  nand g836 (n_859, n_858, n_796);
  nand g837 (n_860, n_855, n_800);
  nand g838 (n_2079, n_859, n_860);
  xor g839 (n_861, B[13], A[20]);
  nand g840 (n_862, n_861, n_796);
  nand g841 (n_863, n_858, n_800);
  nand g842 (n_2117, n_862, n_863);
  xor g843 (n_864, B[13], A[21]);
  nand g844 (n_865, n_864, n_796);
  nand g845 (n_866, n_861, n_800);
  nand g846 (n_2144, n_865, n_866);
  xor g847 (n_867, B[13], A[22]);
  nand g848 (n_868, n_867, n_796);
  nand g849 (n_869, n_864, n_800);
  nand g850 (n_2178, n_868, n_869);
  xor g851 (n_870, B[13], A[23]);
  nand g852 (n_871, n_870, n_796);
  nand g853 (n_872, n_867, n_800);
  nand g854 (n_2203, n_871, n_872);
  xor g855 (n_873, B[13], A[24]);
  nand g856 (n_874, n_873, n_796);
  nand g857 (n_875, n_870, n_800);
  nand g858 (n_2232, n_874, n_875);
  xor g859 (n_876, B[13], A[25]);
  nand g860 (n_877, n_876, n_796);
  nand g861 (n_878, n_873, n_800);
  nand g862 (n_2255, n_877, n_878);
  nand g864 (n_881, B[13], n_796);
  nand g865 (n_882, n_876, n_800);
  nand g866 (n_2277, n_881, n_882);
  nand g869 (n_886, B[13], n_800);
  nand g870 (n_887, n_881, n_886);
  or g874 (n_892, n_890, n_891);
  and g875 (n_1649, B[13], n_892);
  xor g876 (n_893, B[14], B[13]);
  xor g877 (n_895, B[15], B[14]);
  nor g881 (n_988, B[13], B[14]);
  nand g882 (n_986, B[13], B[14]);
  xor g888 (n_901, B[15], A[1]);
  xor g892 (n_904, B[15], A[2]);
  nand g893 (n_905, n_904, n_893);
  nand g894 (n_906, n_901, n_897);
  nand g895 (n_1681, n_905, n_906);
  xor g896 (n_907, B[15], A[3]);
  nand g897 (n_908, n_907, n_893);
  nand g898 (n_909, n_904, n_897);
  nand g899 (n_1694, n_908, n_909);
  xor g900 (n_910, B[15], A[4]);
  nand g901 (n_911, n_910, n_893);
  nand g902 (n_912, n_907, n_897);
  nand g903 (n_1717, n_911, n_912);
  xor g904 (n_913, B[15], A[5]);
  nand g905 (n_914, n_913, n_893);
  nand g906 (n_915, n_910, n_897);
  nand g907 (n_1733, n_914, n_915);
  xor g908 (n_916, B[15], A[6]);
  nand g909 (n_917, n_916, n_893);
  nand g910 (n_918, n_913, n_897);
  nand g911 (n_1755, n_917, n_918);
  xor g912 (n_919, B[15], A[7]);
  nand g913 (n_920, n_919, n_893);
  nand g914 (n_921, n_916, n_897);
  nand g915 (n_1782, n_920, n_921);
  xor g916 (n_922, B[15], A[8]);
  nand g917 (n_923, n_922, n_893);
  nand g918 (n_924, n_919, n_897);
  nand g919 (n_1801, n_923, n_924);
  xor g920 (n_925, B[15], A[9]);
  nand g921 (n_926, n_925, n_893);
  nand g922 (n_927, n_922, n_897);
  nand g923 (n_1829, n_926, n_927);
  xor g924 (n_928, B[15], A[10]);
  nand g925 (n_929, n_928, n_893);
  nand g926 (n_930, n_925, n_897);
  nand g927 (n_1857, n_929, n_930);
  xor g928 (n_931, B[15], A[11]);
  nand g929 (n_932, n_931, n_893);
  nand g930 (n_933, n_928, n_897);
  nand g931 (n_1879, n_932, n_933);
  xor g932 (n_934, B[15], A[12]);
  nand g933 (n_935, n_934, n_893);
  nand g934 (n_936, n_931, n_897);
  nand g935 (n_1913, n_935, n_936);
  xor g936 (n_937, B[15], A[13]);
  nand g937 (n_938, n_937, n_893);
  nand g938 (n_939, n_934, n_897);
  nand g939 (n_1940, n_938, n_939);
  xor g940 (n_940, B[15], A[14]);
  nand g941 (n_941, n_940, n_893);
  nand g942 (n_942, n_937, n_897);
  nand g943 (n_1978, n_941, n_942);
  xor g944 (n_943, B[15], A[15]);
  nand g945 (n_944, n_943, n_893);
  nand g946 (n_945, n_940, n_897);
  nand g947 (n_2007, n_944, n_945);
  xor g948 (n_946, B[15], A[16]);
  nand g949 (n_947, n_946, n_893);
  nand g950 (n_948, n_943, n_897);
  nand g951 (n_2043, n_947, n_948);
  xor g952 (n_949, B[15], A[17]);
  nand g953 (n_950, n_949, n_893);
  nand g954 (n_951, n_946, n_897);
  nand g955 (n_2075, n_950, n_951);
  xor g956 (n_952, B[15], A[18]);
  nand g957 (n_953, n_952, n_893);
  nand g958 (n_954, n_949, n_897);
  nand g959 (n_2111, n_953, n_954);
  xor g960 (n_955, B[15], A[19]);
  nand g961 (n_956, n_955, n_893);
  nand g962 (n_957, n_952, n_897);
  nand g963 (n_2140, n_956, n_957);
  xor g964 (n_958, B[15], A[20]);
  nand g965 (n_959, n_958, n_893);
  nand g966 (n_960, n_955, n_897);
  nand g967 (n_2172, n_959, n_960);
  xor g968 (n_961, B[15], A[21]);
  nand g969 (n_962, n_961, n_893);
  nand g970 (n_963, n_958, n_897);
  nand g971 (n_2200, n_962, n_963);
  xor g972 (n_964, B[15], A[22]);
  nand g973 (n_965, n_964, n_893);
  nand g974 (n_966, n_961, n_897);
  nand g975 (n_2230, n_965, n_966);
  xor g976 (n_967, B[15], A[23]);
  nand g977 (n_968, n_967, n_893);
  nand g978 (n_969, n_964, n_897);
  nand g979 (n_2253, n_968, n_969);
  xor g980 (n_970, B[15], A[24]);
  nand g981 (n_971, n_970, n_893);
  nand g982 (n_972, n_967, n_897);
  nand g983 (n_2279, n_971, n_972);
  xor g984 (n_973, B[15], A[25]);
  nand g985 (n_974, n_973, n_893);
  nand g986 (n_975, n_970, n_897);
  nand g987 (n_2305, n_974, n_975);
  nand g989 (n_978, B[15], n_893);
  nand g990 (n_979, n_973, n_897);
  nand g991 (n_2324, n_978, n_979);
  nand g994 (n_983, B[15], n_897);
  nand g995 (n_984, n_978, n_983);
  or g999 (n_989, n_987, n_988);
  and g1000 (n_1677, B[15], n_989);
  xor g1001 (n_990, B[16], B[15]);
  xor g1002 (n_992, B[17], B[16]);
  nor g1006 (n_1085, B[15], B[16]);
  nand g1007 (n_1083, B[15], B[16]);
  xor g1013 (n_998, B[17], A[1]);
  xor g1017 (n_1001, B[17], A[2]);
  nand g1018 (n_1002, n_1001, n_990);
  nand g1019 (n_1003, n_998, n_994);
  nand g1020 (n_1718, n_1002, n_1003);
  xor g1021 (n_1004, B[17], A[3]);
  nand g1022 (n_1005, n_1004, n_990);
  nand g1023 (n_1006, n_1001, n_994);
  nand g1024 (n_1731, n_1005, n_1006);
  xor g1025 (n_1007, B[17], A[4]);
  nand g1026 (n_1008, n_1007, n_990);
  nand g1027 (n_1009, n_1004, n_994);
  nand g1028 (n_1753, n_1008, n_1009);
  xor g1029 (n_1010, B[17], A[5]);
  nand g1030 (n_1011, n_1010, n_990);
  nand g1031 (n_1012, n_1007, n_994);
  nand g1032 (n_1776, n_1011, n_1012);
  xor g1033 (n_1013, B[17], A[6]);
  nand g1034 (n_1014, n_1013, n_990);
  nand g1035 (n_1015, n_1010, n_994);
  nand g1036 (n_1802, n_1014, n_1015);
  xor g1037 (n_1016, B[17], A[7]);
  nand g1038 (n_1017, n_1016, n_990);
  nand g1039 (n_1018, n_1013, n_994);
  nand g1040 (n_1832, n_1017, n_1018);
  xor g1041 (n_1019, B[17], A[8]);
  nand g1042 (n_1020, n_1019, n_990);
  nand g1043 (n_1021, n_1016, n_994);
  nand g1044 (n_1853, n_1020, n_1021);
  xor g1045 (n_1022, B[17], A[9]);
  nand g1046 (n_1023, n_1022, n_990);
  nand g1047 (n_1024, n_1019, n_994);
  nand g1048 (n_1885, n_1023, n_1024);
  xor g1049 (n_1025, B[17], A[10]);
  nand g1050 (n_1026, n_1025, n_990);
  nand g1051 (n_1027, n_1022, n_994);
  nand g1052 (n_1918, n_1026, n_1027);
  xor g1053 (n_1028, B[17], A[11]);
  nand g1054 (n_1029, n_1028, n_990);
  nand g1055 (n_1030, n_1025, n_994);
  nand g1056 (n_1947, n_1029, n_1030);
  xor g1057 (n_1031, B[17], A[12]);
  nand g1058 (n_1032, n_1031, n_990);
  nand g1059 (n_1033, n_1028, n_994);
  nand g1060 (n_1979, n_1032, n_1033);
  xor g1061 (n_1034, B[17], A[13]);
  nand g1062 (n_1035, n_1034, n_990);
  nand g1063 (n_1036, n_1031, n_994);
  nand g1064 (n_2016, n_1035, n_1036);
  xor g1065 (n_1037, B[17], A[14]);
  nand g1066 (n_1038, n_1037, n_990);
  nand g1067 (n_1039, n_1034, n_994);
  nand g1068 (n_2049, n_1038, n_1039);
  xor g1069 (n_1040, B[17], A[15]);
  nand g1070 (n_1041, n_1040, n_990);
  nand g1071 (n_1042, n_1037, n_994);
  nand g1072 (n_2084, n_1041, n_1042);
  xor g1073 (n_1043, B[17], A[16]);
  nand g1074 (n_1044, n_1043, n_990);
  nand g1075 (n_1045, n_1040, n_994);
  nand g1076 (n_2118, n_1044, n_1045);
  xor g1077 (n_1046, B[17], A[17]);
  nand g1078 (n_1047, n_1046, n_990);
  nand g1079 (n_1048, n_1043, n_994);
  nand g1080 (n_2146, n_1047, n_1048);
  xor g1081 (n_1049, B[17], A[18]);
  nand g1082 (n_1050, n_1049, n_990);
  nand g1083 (n_1051, n_1046, n_994);
  nand g1084 (n_2173, n_1050, n_1051);
  xor g1085 (n_1052, B[17], A[19]);
  nand g1086 (n_1053, n_1052, n_990);
  nand g1087 (n_1054, n_1049, n_994);
  nand g1088 (n_2199, n_1053, n_1054);
  xor g1089 (n_1055, B[17], A[20]);
  nand g1090 (n_1056, n_1055, n_990);
  nand g1091 (n_1057, n_1052, n_994);
  nand g1092 (n_2234, n_1056, n_1057);
  xor g1093 (n_1058, B[17], A[21]);
  nand g1094 (n_1059, n_1058, n_990);
  nand g1095 (n_1060, n_1055, n_994);
  nand g1096 (n_2252, n_1059, n_1060);
  xor g1097 (n_1061, B[17], A[22]);
  nand g1098 (n_1062, n_1061, n_990);
  nand g1099 (n_1063, n_1058, n_994);
  nand g1100 (n_2281, n_1062, n_1063);
  xor g1101 (n_1064, B[17], A[23]);
  nand g1102 (n_1065, n_1064, n_990);
  nand g1103 (n_1066, n_1061, n_994);
  nand g1104 (n_2301, n_1065, n_1066);
  xor g1105 (n_1067, B[17], A[24]);
  nand g1106 (n_1068, n_1067, n_990);
  nand g1107 (n_1069, n_1064, n_994);
  nand g1108 (n_2325, n_1068, n_1069);
  xor g1109 (n_1070, B[17], A[25]);
  nand g1110 (n_1071, n_1070, n_990);
  nand g1111 (n_1072, n_1067, n_994);
  nand g1112 (n_2345, n_1071, n_1072);
  nand g1114 (n_1075, B[17], n_990);
  nand g1115 (n_1076, n_1070, n_994);
  nand g1116 (n_2361, n_1075, n_1076);
  nand g1119 (n_1080, B[17], n_994);
  nand g1120 (n_1081, n_1075, n_1080);
  or g1124 (n_1086, n_1084, n_1085);
  and g1125 (n_1711, B[17], n_1086);
  xor g1126 (n_1087, B[18], B[17]);
  xor g1127 (n_1089, B[19], B[18]);
  nor g1131 (n_1182, B[17], B[18]);
  nand g1132 (n_1180, B[17], B[18]);
  xor g1138 (n_1095, B[19], A[1]);
  xor g1142 (n_1098, B[19], A[2]);
  nand g1143 (n_1099, n_1098, n_1087);
  nand g1144 (n_1100, n_1095, n_1091);
  nand g1145 (n_1760, n_1099, n_1100);
  xor g1146 (n_1101, B[19], A[3]);
  nand g1147 (n_1102, n_1101, n_1087);
  nand g1148 (n_1103, n_1098, n_1091);
  nand g1149 (n_1774, n_1102, n_1103);
  xor g1150 (n_1104, B[19], A[4]);
  nand g1151 (n_1105, n_1104, n_1087);
  nand g1152 (n_1106, n_1101, n_1091);
  nand g1153 (n_1799, n_1105, n_1106);
  xor g1154 (n_1107, B[19], A[5]);
  nand g1155 (n_1108, n_1107, n_1087);
  nand g1156 (n_1109, n_1104, n_1091);
  nand g1157 (n_1825, n_1108, n_1109);
  xor g1158 (n_1110, B[19], A[6]);
  nand g1159 (n_1111, n_1110, n_1087);
  nand g1160 (n_1112, n_1107, n_1091);
  nand g1161 (n_1852, n_1111, n_1112);
  xor g1162 (n_1113, B[19], A[7]);
  nand g1163 (n_1114, n_1113, n_1087);
  nand g1164 (n_1115, n_1110, n_1091);
  nand g1165 (n_1888, n_1114, n_1115);
  xor g1166 (n_1116, B[19], A[8]);
  nand g1167 (n_1117, n_1116, n_1087);
  nand g1168 (n_1118, n_1113, n_1091);
  nand g1169 (n_1911, n_1117, n_1118);
  xor g1170 (n_1119, B[19], A[9]);
  nand g1171 (n_1120, n_1119, n_1087);
  nand g1172 (n_1121, n_1116, n_1091);
  nand g1173 (n_1939, n_1120, n_1121);
  xor g1174 (n_1122, B[19], A[10]);
  nand g1175 (n_1123, n_1122, n_1087);
  nand g1176 (n_1124, n_1119, n_1091);
  nand g1177 (n_1981, n_1123, n_1124);
  xor g1178 (n_1125, B[19], A[11]);
  nand g1179 (n_1126, n_1125, n_1087);
  nand g1180 (n_1127, n_1122, n_1091);
  nand g1181 (n_2011, n_1126, n_1127);
  xor g1182 (n_1128, B[19], A[12]);
  nand g1183 (n_1129, n_1128, n_1087);
  nand g1184 (n_1130, n_1125, n_1091);
  nand g1185 (n_2048, n_1129, n_1130);
  xor g1186 (n_1131, B[19], A[13]);
  nand g1187 (n_1132, n_1131, n_1087);
  nand g1188 (n_1133, n_1128, n_1091);
  nand g1189 (n_2080, n_1132, n_1133);
  xor g1190 (n_1134, B[19], A[14]);
  nand g1191 (n_1135, n_1134, n_1087);
  nand g1192 (n_1136, n_1131, n_1091);
  nand g1193 (n_2109, n_1135, n_1136);
  xor g1194 (n_1137, B[19], A[15]);
  nand g1195 (n_1138, n_1137, n_1087);
  nand g1196 (n_1139, n_1134, n_1091);
  nand g1197 (n_2145, n_1138, n_1139);
  xor g1198 (n_1140, B[19], A[16]);
  nand g1199 (n_1141, n_1140, n_1087);
  nand g1200 (n_1142, n_1137, n_1091);
  nand g1201 (n_2171, n_1141, n_1142);
  xor g1202 (n_1143, B[19], A[17]);
  nand g1203 (n_1144, n_1143, n_1087);
  nand g1204 (n_1145, n_1140, n_1091);
  nand g1205 (n_2202, n_1144, n_1145);
  xor g1206 (n_1146, B[19], A[18]);
  nand g1207 (n_1147, n_1146, n_1087);
  nand g1208 (n_1148, n_1143, n_1091);
  nand g1209 (n_2233, n_1147, n_1148);
  xor g1210 (n_1149, B[19], A[19]);
  nand g1211 (n_1150, n_1149, n_1087);
  nand g1212 (n_1151, n_1146, n_1091);
  nand g1213 (n_2254, n_1150, n_1151);
  xor g1214 (n_1152, B[19], A[20]);
  nand g1215 (n_1153, n_1152, n_1087);
  nand g1216 (n_1154, n_1149, n_1091);
  nand g1217 (n_2282, n_1153, n_1154);
  xor g1218 (n_1155, B[19], A[21]);
  nand g1219 (n_1156, n_1155, n_1087);
  nand g1220 (n_1157, n_1152, n_1091);
  nand g1221 (n_2299, n_1156, n_1157);
  xor g1222 (n_1158, B[19], A[22]);
  nand g1223 (n_1159, n_1158, n_1087);
  nand g1224 (n_1160, n_1155, n_1091);
  nand g1225 (n_2323, n_1159, n_1160);
  xor g1226 (n_1161, B[19], A[23]);
  nand g1227 (n_1162, n_1161, n_1087);
  nand g1228 (n_1163, n_1158, n_1091);
  nand g1229 (n_2340, n_1162, n_1163);
  xor g1230 (n_1164, B[19], A[24]);
  nand g1231 (n_1165, n_1164, n_1087);
  nand g1232 (n_1166, n_1161, n_1091);
  nand g1233 (n_2362, n_1165, n_1166);
  xor g1234 (n_1167, B[19], A[25]);
  nand g1235 (n_1168, n_1167, n_1087);
  nand g1236 (n_1169, n_1164, n_1091);
  nand g1237 (n_2379, n_1168, n_1169);
  nand g1239 (n_1172, B[19], n_1087);
  nand g1240 (n_1173, n_1167, n_1091);
  nand g1241 (n_2391, n_1172, n_1173);
  nand g1244 (n_1177, B[19], n_1091);
  nand g1245 (n_1178, n_1172, n_1177);
  or g1249 (n_1183, n_1181, n_1182);
  and g1250 (n_1751, B[19], n_1183);
  xor g1251 (n_1184, B[20], B[19]);
  xor g1252 (n_1186, B[21], B[20]);
  nor g1256 (n_1279, B[19], B[20]);
  nand g1257 (n_1277, B[19], B[20]);
  xor g1263 (n_1192, B[21], A[1]);
  xor g1267 (n_1195, B[21], A[2]);
  nand g1268 (n_1196, n_1195, n_1184);
  nand g1269 (n_1197, n_1192, n_1188);
  nand g1270 (n_1807, n_1196, n_1197);
  xor g1271 (n_1198, B[21], A[3]);
  nand g1272 (n_1199, n_1198, n_1184);
  nand g1273 (n_1200, n_1195, n_1188);
  nand g1274 (n_1823, n_1199, n_1200);
  xor g1275 (n_1201, B[21], A[4]);
  nand g1276 (n_1202, n_1201, n_1184);
  nand g1277 (n_1203, n_1198, n_1188);
  nand g1278 (n_1851, n_1202, n_1203);
  xor g1279 (n_1204, B[21], A[5]);
  nand g1280 (n_1205, n_1204, n_1184);
  nand g1281 (n_1206, n_1201, n_1188);
  nand g1282 (n_1880, n_1205, n_1206);
  xor g1283 (n_1207, B[21], A[6]);
  nand g1284 (n_1208, n_1207, n_1184);
  nand g1285 (n_1209, n_1204, n_1188);
  nand g1286 (n_1910, n_1208, n_1209);
  xor g1287 (n_1210, B[21], A[7]);
  nand g1288 (n_1211, n_1210, n_1184);
  nand g1289 (n_1212, n_1207, n_1188);
  nand g1290 (n_1946, n_1211, n_1212);
  xor g1291 (n_1213, B[21], A[8]);
  nand g1292 (n_1214, n_1213, n_1184);
  nand g1293 (n_1215, n_1210, n_1188);
  nand g1294 (n_1975, n_1214, n_1215);
  xor g1295 (n_1216, B[21], A[9]);
  nand g1296 (n_1217, n_1216, n_1184);
  nand g1297 (n_1218, n_1213, n_1188);
  nand g1298 (n_2015, n_1217, n_1218);
  xor g1299 (n_1219, B[21], A[10]);
  nand g1300 (n_1220, n_1219, n_1184);
  nand g1301 (n_1221, n_1216, n_1188);
  nand g1302 (n_2044, n_1220, n_1221);
  xor g1303 (n_1222, B[21], A[11]);
  nand g1304 (n_1223, n_1222, n_1184);
  nand g1305 (n_1224, n_1219, n_1188);
  nand g1306 (n_2083, n_1223, n_1224);
  xor g1307 (n_1225, B[21], A[12]);
  nand g1308 (n_1226, n_1225, n_1184);
  nand g1309 (n_1227, n_1222, n_1188);
  nand g1310 (n_2112, n_1226, n_1227);
  xor g1311 (n_1228, B[21], A[13]);
  nand g1312 (n_1229, n_1228, n_1184);
  nand g1313 (n_1230, n_1225, n_1188);
  nand g1314 (n_2148, n_1229, n_1230);
  xor g1315 (n_1231, B[21], A[14]);
  nand g1316 (n_1232, n_1231, n_1184);
  nand g1317 (n_1233, n_1228, n_1188);
  nand g1318 (n_2174, n_1232, n_1233);
  xor g1319 (n_1234, B[21], A[15]);
  nand g1320 (n_1235, n_1234, n_1184);
  nand g1321 (n_1236, n_1231, n_1188);
  nand g1322 (n_2206, n_1235, n_1236);
  xor g1323 (n_1237, B[21], A[16]);
  nand g1324 (n_1238, n_1237, n_1184);
  nand g1325 (n_1239, n_1234, n_1188);
  nand g1326 (n_2229, n_1238, n_1239);
  xor g1327 (n_1240, B[21], A[17]);
  nand g1328 (n_1241, n_1240, n_1184);
  nand g1329 (n_1242, n_1237, n_1188);
  nand g1330 (n_2258, n_1241, n_1242);
  xor g1331 (n_1243, B[21], A[18]);
  nand g1332 (n_1244, n_1243, n_1184);
  nand g1333 (n_1245, n_1240, n_1188);
  nand g1334 (n_2283, n_1244, n_1245);
  xor g1335 (n_1246, B[21], A[19]);
  nand g1336 (n_1247, n_1246, n_1184);
  nand g1337 (n_1248, n_1243, n_1188);
  nand g1338 (n_2302, n_1247, n_1248);
  xor g1339 (n_1249, B[21], A[20]);
  nand g1340 (n_1250, n_1249, n_1184);
  nand g1341 (n_1251, n_1246, n_1188);
  nand g1342 (n_2326, n_1250, n_1251);
  xor g1343 (n_1252, B[21], A[21]);
  nand g1344 (n_1253, n_1252, n_1184);
  nand g1345 (n_1254, n_1249, n_1188);
  nand g1346 (n_2341, n_1253, n_1254);
  xor g1347 (n_1255, B[21], A[22]);
  nand g1348 (n_1256, n_1255, n_1184);
  nand g1349 (n_1257, n_1252, n_1188);
  nand g1350 (n_2360, n_1256, n_1257);
  xor g1351 (n_1258, B[21], A[23]);
  nand g1352 (n_1259, n_1258, n_1184);
  nand g1353 (n_1260, n_1255, n_1188);
  nand g1354 (n_2375, n_1259, n_1260);
  xor g1355 (n_1261, B[21], A[24]);
  nand g1356 (n_1262, n_1261, n_1184);
  nand g1357 (n_1263, n_1258, n_1188);
  nand g1358 (n_2392, n_1262, n_1263);
  xor g1359 (n_1264, B[21], A[25]);
  nand g1360 (n_1265, n_1264, n_1184);
  nand g1361 (n_1266, n_1261, n_1188);
  nand g1362 (n_2404, n_1265, n_1266);
  nand g1364 (n_1269, B[21], n_1184);
  nand g1365 (n_1270, n_1264, n_1188);
  nand g1366 (n_2419, n_1269, n_1270);
  nand g1369 (n_1274, B[21], n_1188);
  nand g1370 (n_1275, n_1269, n_1274);
  or g1374 (n_1280, n_1278, n_1279);
  and g1375 (n_1797, B[21], n_1280);
  xor g1376 (n_1281, B[22], B[21]);
  xor g1377 (n_1283, B[23], B[22]);
  nor g1381 (n_1376, B[21], B[22]);
  nand g1382 (n_1374, B[21], B[22]);
  xor g1388 (n_1289, B[23], A[1]);
  xor g1392 (n_1292, B[23], A[2]);
  nand g1393 (n_1293, n_1292, n_1281);
  nand g1394 (n_1294, n_1289, n_1285);
  nand g1395 (n_1860, n_1293, n_1294);
  xor g1396 (n_1295, B[23], A[3]);
  nand g1397 (n_1296, n_1295, n_1281);
  nand g1398 (n_1297, n_1292, n_1285);
  nand g1399 (n_1878, n_1296, n_1297);
  xor g1400 (n_1298, B[23], A[4]);
  nand g1401 (n_1299, n_1298, n_1281);
  nand g1402 (n_1300, n_1295, n_1285);
  nand g1403 (n_1909, n_1299, n_1300);
  xor g1404 (n_1301, B[23], A[5]);
  nand g1405 (n_1302, n_1301, n_1281);
  nand g1406 (n_1303, n_1298, n_1285);
  nand g1407 (n_1950, n_1302, n_1303);
  xor g1408 (n_1304, B[23], A[6]);
  nand g1409 (n_1305, n_1304, n_1281);
  nand g1410 (n_1306, n_1301, n_1285);
  nand g1411 (n_1976, n_1305, n_1306);
  xor g1412 (n_1307, B[23], A[7]);
  nand g1413 (n_1308, n_1307, n_1281);
  nand g1414 (n_1309, n_1304, n_1285);
  nand g1415 (n_2014, n_1308, n_1309);
  xor g1416 (n_1310, B[23], A[8]);
  nand g1417 (n_1311, n_1310, n_1281);
  nand g1418 (n_1312, n_1307, n_1285);
  nand g1419 (n_2045, n_1311, n_1312);
  xor g1420 (n_1313, B[23], A[9]);
  nand g1421 (n_1314, n_1313, n_1281);
  nand g1422 (n_1315, n_1310, n_1285);
  nand g1423 (n_2082, n_1314, n_1315);
  xor g1424 (n_1316, B[23], A[10]);
  nand g1425 (n_1317, n_1316, n_1281);
  nand g1426 (n_1318, n_1313, n_1285);
  nand g1427 (n_2115, n_1317, n_1318);
  xor g1428 (n_1319, B[23], A[11]);
  nand g1429 (n_1320, n_1319, n_1281);
  nand g1430 (n_1321, n_1316, n_1285);
  nand g1431 (n_2147, n_1320, n_1321);
  xor g1432 (n_1322, B[23], A[12]);
  nand g1433 (n_1323, n_1322, n_1281);
  nand g1434 (n_1324, n_1319, n_1285);
  nand g1435 (n_2176, n_1323, n_1324);
  xor g1436 (n_1325, B[23], A[13]);
  nand g1437 (n_1326, n_1325, n_1281);
  nand g1438 (n_1327, n_1322, n_1285);
  nand g1439 (n_2205, n_1326, n_1327);
  xor g1440 (n_1328, B[23], A[14]);
  nand g1441 (n_1329, n_1328, n_1281);
  nand g1442 (n_1330, n_1325, n_1285);
  nand g1443 (n_2231, n_1329, n_1330);
  xor g1444 (n_1331, B[23], A[15]);
  nand g1445 (n_1332, n_1331, n_1281);
  nand g1446 (n_1333, n_1328, n_1285);
  nand g1447 (n_2257, n_1332, n_1333);
  xor g1448 (n_1334, B[23], A[16]);
  nand g1449 (n_1335, n_1334, n_1281);
  nand g1450 (n_1336, n_1331, n_1285);
  nand g1451 (n_2280, n_1335, n_1336);
  xor g1452 (n_1337, B[23], A[17]);
  nand g1453 (n_1338, n_1337, n_1281);
  nand g1454 (n_1339, n_1334, n_1285);
  nand g1455 (n_2303, n_1338, n_1339);
  xor g1456 (n_1340, B[23], A[18]);
  nand g1457 (n_1341, n_1340, n_1281);
  nand g1458 (n_1342, n_1337, n_1285);
  nand g1459 (n_2322, n_1341, n_1342);
  xor g1460 (n_1343, B[23], A[19]);
  nand g1461 (n_1344, n_1343, n_1281);
  nand g1462 (n_1345, n_1340, n_1285);
  nand g1463 (n_2343, n_1344, n_1345);
  xor g1464 (n_1346, B[23], A[20]);
  nand g1465 (n_1347, n_1346, n_1281);
  nand g1466 (n_1348, n_1343, n_1285);
  nand g1467 (n_2363, n_1347, n_1348);
  xor g1468 (n_1349, B[23], A[21]);
  nand g1469 (n_1350, n_1349, n_1281);
  nand g1470 (n_1351, n_1346, n_1285);
  nand g1471 (n_2378, n_1350, n_1351);
  xor g1472 (n_1352, B[23], A[22]);
  nand g1473 (n_1353, n_1352, n_1281);
  nand g1474 (n_1354, n_1349, n_1285);
  nand g1475 (n_2394, n_1353, n_1354);
  xor g1476 (n_1355, B[23], A[23]);
  nand g1477 (n_1356, n_1355, n_1281);
  nand g1478 (n_1357, n_1352, n_1285);
  nand g1479 (n_2407, n_1356, n_1357);
  xor g1480 (n_1358, B[23], A[24]);
  nand g1481 (n_1359, n_1358, n_1281);
  nand g1482 (n_1360, n_1355, n_1285);
  nand g1483 (n_2417, n_1359, n_1360);
  xor g1484 (n_1361, B[23], A[25]);
  nand g1485 (n_1362, n_1361, n_1281);
  nand g1486 (n_1363, n_1358, n_1285);
  nand g1487 (n_2427, n_1362, n_1363);
  nand g1489 (n_1366, B[23], n_1281);
  nand g1490 (n_1367, n_1361, n_1285);
  nand g1491 (n_2438, n_1366, n_1367);
  nand g1494 (n_1371, B[23], n_1285);
  nand g1495 (n_1372, n_1366, n_1371);
  or g1499 (n_1377, n_1375, n_1376);
  and g1500 (n_1849, B[23], n_1377);
  xor g1501 (n_1378, B[24], B[23]);
  xor g1502 (n_1380, B[25], B[24]);
  nor g1506 (n_1473, B[23], B[24]);
  nand g1507 (n_1471, B[23], B[24]);
  xor g1513 (n_1386, B[25], A[1]);
  xor g1517 (n_1389, B[25], A[2]);
  nand g1518 (n_1390, n_1389, n_1378);
  nand g1519 (n_1391, n_1386, n_1382);
  nand g1520 (n_1919, n_1390, n_1391);
  xor g1521 (n_1392, B[25], A[3]);
  nand g1522 (n_1393, n_1392, n_1378);
  nand g1523 (n_1394, n_1389, n_1382);
  nand g1524 (n_1941, n_1393, n_1394);
  xor g1525 (n_1395, B[25], A[4]);
  nand g1526 (n_1396, n_1395, n_1378);
  nand g1527 (n_1397, n_1392, n_1382);
  nand g1528 (n_1972, n_1396, n_1397);
  xor g1529 (n_1398, B[25], A[5]);
  nand g1530 (n_1399, n_1398, n_1378);
  nand g1531 (n_1400, n_1395, n_1382);
  nand g1532 (n_2009, n_1399, n_1400);
  xor g1533 (n_1401, B[25], A[6]);
  nand g1534 (n_1402, n_1401, n_1378);
  nand g1535 (n_1403, n_1398, n_1382);
  nand g1536 (n_2041, n_1402, n_1403);
  xor g1537 (n_1404, B[25], A[7]);
  nand g1538 (n_1405, n_1404, n_1378);
  nand g1539 (n_1406, n_1401, n_1382);
  nand g1540 (n_2078, n_1405, n_1406);
  xor g1541 (n_1407, B[25], A[8]);
  nand g1542 (n_1408, n_1407, n_1378);
  nand g1543 (n_1409, n_1404, n_1382);
  nand g1544 (n_2113, n_1408, n_1409);
  xor g1545 (n_1410, B[25], A[9]);
  nand g1546 (n_1411, n_1410, n_1378);
  nand g1547 (n_1412, n_1407, n_1382);
  nand g1548 (n_2143, n_1411, n_1412);
  xor g1549 (n_1413, B[25], A[10]);
  nand g1550 (n_1414, n_1413, n_1378);
  nand g1551 (n_1415, n_1410, n_1382);
  nand g1552 (n_2175, n_1414, n_1415);
  xor g1553 (n_1416, B[25], A[11]);
  nand g1554 (n_1417, n_1416, n_1378);
  nand g1555 (n_1418, n_1413, n_1382);
  nand g1556 (n_2201, n_1417, n_1418);
  xor g1557 (n_1419, B[25], A[12]);
  nand g1558 (n_1420, n_1419, n_1378);
  nand g1559 (n_1421, n_1416, n_1382);
  nand g1560 (n_2228, n_1420, n_1421);
  xor g1561 (n_1422, B[25], A[13]);
  nand g1562 (n_1423, n_1422, n_1378);
  nand g1563 (n_1424, n_1419, n_1382);
  nand g1564 (n_2259, n_1423, n_1424);
  xor g1565 (n_1425, B[25], A[14]);
  nand g1566 (n_1426, n_1425, n_1378);
  nand g1567 (n_1427, n_1422, n_1382);
  nand g1568 (n_2278, n_1426, n_1427);
  xor g1569 (n_1428, B[25], A[15]);
  nand g1570 (n_1429, n_1428, n_1378);
  nand g1571 (n_1430, n_1425, n_1382);
  nand g1572 (n_2304, n_1429, n_1430);
  xor g1573 (n_1431, B[25], A[16]);
  nand g1574 (n_1432, n_1431, n_1378);
  nand g1575 (n_1433, n_1428, n_1382);
  nand g1576 (n_2321, n_1432, n_1433);
  xor g1577 (n_1434, B[25], A[17]);
  nand g1578 (n_1435, n_1434, n_1378);
  nand g1579 (n_1436, n_1431, n_1382);
  nand g1580 (n_2342, n_1435, n_1436);
  xor g1581 (n_1437, B[25], A[18]);
  nand g1582 (n_1438, n_1437, n_1378);
  nand g1583 (n_1439, n_1434, n_1382);
  nand g1584 (n_2359, n_1438, n_1439);
  xor g1585 (n_1440, B[25], A[19]);
  nand g1586 (n_1441, n_1440, n_1378);
  nand g1587 (n_1442, n_1437, n_1382);
  nand g1588 (n_2377, n_1441, n_1442);
  xor g1589 (n_1443, B[25], A[20]);
  nand g1590 (n_1444, n_1443, n_1378);
  nand g1591 (n_1445, n_1440, n_1382);
  nand g1592 (n_2393, n_1444, n_1445);
  xor g1593 (n_1446, B[25], A[21]);
  nand g1594 (n_1447, n_1446, n_1378);
  nand g1595 (n_1448, n_1443, n_1382);
  nand g1596 (n_2406, n_1447, n_1448);
  xor g1597 (n_1449, B[25], A[22]);
  nand g1598 (n_1450, n_1449, n_1378);
  nand g1599 (n_1451, n_1446, n_1382);
  nand g1600 (n_2418, n_1450, n_1451);
  xor g1601 (n_1452, B[25], A[23]);
  nand g1602 (n_1453, n_1452, n_1378);
  nand g1603 (n_1454, n_1449, n_1382);
  nand g1604 (n_2428, n_1453, n_1454);
  xor g1605 (n_1455, B[25], A[24]);
  nand g1606 (n_1456, n_1455, n_1378);
  nand g1607 (n_1457, n_1452, n_1382);
  nand g1608 (n_2437, n_1456, n_1457);
  xor g1609 (n_1458, B[25], A[25]);
  nand g1610 (n_1459, n_1458, n_1378);
  nand g1611 (n_1460, n_1455, n_1382);
  nand g1612 (n_2445, n_1459, n_1460);
  nand g1614 (n_1463, B[25], n_1378);
  nand g1615 (n_1464, n_1458, n_1382);
  nand g1616 (n_2451, n_1463, n_1464);
  nand g1619 (n_1468, B[25], n_1382);
  nand g1620 (n_1469, n_1463, n_1468);
  or g1624 (n_1474, n_1472, n_1473);
  and g1625 (n_1907, B[25], n_1474);
  nand g1643 (n_1497, A[2], B[25]);
  nand g1647 (n_1501, A[3], B[25]);
  nand g1651 (n_1505, A[4], B[25]);
  nand g1655 (n_1509, A[5], B[25]);
  nand g1659 (n_1513, A[6], B[25]);
  nand g1663 (n_1517, A[7], B[25]);
  nand g1667 (n_1521, A[8], B[25]);
  nand g1671 (n_1525, A[9], B[25]);
  nand g1675 (n_1529, A[10], B[25]);
  nand g1679 (n_1533, A[11], B[25]);
  nand g1683 (n_1537, A[12], B[25]);
  nand g1687 (n_1541, A[13], B[25]);
  nand g1691 (n_1545, A[14], B[25]);
  nand g1695 (n_1549, A[15], B[25]);
  nand g1699 (n_1553, A[16], B[25]);
  nand g1703 (n_1557, A[17], B[25]);
  nand g1707 (n_1561, A[18], B[25]);
  nand g1711 (n_1565, A[19], B[25]);
  nand g1715 (n_1569, A[20], B[25]);
  nand g1719 (n_1573, A[21], B[25]);
  nand g1723 (n_1577, A[22], B[25]);
  nand g1727 (n_1581, A[23], B[25]);
  nand g1731 (n_1585, A[24], B[25]);
  xor g2040 (n_202, n_1597, n_1598);
  and g2041 (n_149, n_1597, n_1598);
  xor g2042 (n_201, n_1599, n_1600);
  and g2043 (n_148, n_1599, n_1600);
  xor g2044 (n_1605, n_1601, n_1602);
  and g2045 (n_1610, n_1601, n_1602);
  xor g2046 (n_2457, n_1603, n_1604);
  xor g2047 (n_200, n_2457, n_1605);
  nand g2048 (n_2458, n_1603, n_1604);
  nand g2049 (n_2459, n_1605, n_1604);
  nand g2050 (n_2460, n_1603, n_1605);
  nand g2051 (n_147, n_2458, n_2459, n_2460);
  xor g2052 (n_1609, n_1606, n_1607);
  and g2053 (n_1617, n_1606, n_1607);
  xor g2054 (n_2461, n_1608, n_1609);
  xor g2055 (n_199, n_2461, n_1610);
  nand g2056 (n_2462, n_1608, n_1609);
  nand g2057 (n_2463, n_1610, n_1609);
  nand g2058 (n_2464, n_1608, n_1610);
  nand g2059 (n_146, n_2462, n_2463, n_2464);
  xor g2060 (n_1616, n_1611, n_1612);
  and g2061 (n_1623, n_1611, n_1612);
  xor g2062 (n_2465, n_1613, n_1614);
  xor g2063 (n_1618, n_2465, n_1615);
  nand g2064 (n_2466, n_1613, n_1614);
  nand g2065 (n_2467, n_1615, n_1614);
  nand g2066 (n_2468, n_1613, n_1615);
  nand g2067 (n_1625, n_2466, n_2467, n_2468);
  xor g2068 (n_2469, n_1616, n_1617);
  xor g2069 (n_198, n_2469, n_1618);
  nand g2070 (n_2470, n_1616, n_1617);
  nand g2071 (n_2471, n_1618, n_1617);
  nand g2072 (n_2472, n_1616, n_1618);
  nand g2073 (n_145, n_2470, n_2471, n_2472);
  xor g2074 (n_1624, n_1619, n_1620);
  and g2075 (n_1634, n_1619, n_1620);
  xor g2076 (n_2473, n_1621, n_1622);
  xor g2077 (n_1626, n_2473, n_1623);
  nand g2078 (n_2474, n_1621, n_1622);
  nand g2079 (n_2475, n_1623, n_1622);
  nand g2080 (n_2476, n_1621, n_1623);
  nand g2081 (n_1636, n_2474, n_2475, n_2476);
  xor g2082 (n_2477, n_1624, n_1625);
  xor g2083 (n_197, n_2477, n_1626);
  nand g2084 (n_2478, n_1624, n_1625);
  nand g2085 (n_2479, n_1626, n_1625);
  nand g2086 (n_2480, n_1624, n_1626);
  nand g2087 (n_144, n_2478, n_2479, n_2480);
  xor g2088 (n_1633, n_1627, n_1628);
  and g2089 (n_1644, n_1627, n_1628);
  xor g2090 (n_2481, n_1629, n_1630);
  xor g2091 (n_1635, n_2481, n_1631);
  nand g2092 (n_2482, n_1629, n_1630);
  nand g2093 (n_2483, n_1631, n_1630);
  nand g2094 (n_2484, n_1629, n_1631);
  nand g2095 (n_1645, n_2482, n_2483, n_2484);
  xor g2096 (n_2485, n_1632, n_1633);
  xor g2097 (n_1637, n_2485, n_1634);
  nand g2098 (n_2486, n_1632, n_1633);
  nand g2099 (n_2487, n_1634, n_1633);
  nand g2100 (n_2488, n_1632, n_1634);
  nand g2101 (n_1647, n_2486, n_2487, n_2488);
  xor g2102 (n_2489, n_1635, n_1636);
  xor g2103 (n_196, n_2489, n_1637);
  nand g2104 (n_2490, n_1635, n_1636);
  nand g2105 (n_2491, n_1637, n_1636);
  nand g2106 (n_2492, n_1635, n_1637);
  nand g2107 (n_143, n_2490, n_2491, n_2492);
  xor g2108 (n_1643, n_1638, n_1639);
  and g2109 (n_1657, n_1638, n_1639);
  xor g2110 (n_2493, n_1640, n_1641);
  xor g2111 (n_1646, n_2493, n_1642);
  nand g2112 (n_2494, n_1640, n_1641);
  nand g2113 (n_2495, n_1642, n_1641);
  nand g2114 (n_2496, n_1640, n_1642);
  nand g2115 (n_1658, n_2494, n_2495, n_2496);
  xor g2116 (n_2497, n_1643, n_1644);
  xor g2117 (n_1648, n_2497, n_1645);
  nand g2118 (n_2498, n_1643, n_1644);
  nand g2119 (n_2499, n_1645, n_1644);
  nand g2120 (n_2500, n_1643, n_1645);
  nand g2121 (n_1661, n_2498, n_2499, n_2500);
  xor g2122 (n_2501, n_1646, n_1647);
  xor g2123 (n_195, n_2501, n_1648);
  nand g2124 (n_2502, n_1646, n_1647);
  nand g2125 (n_2503, n_1648, n_1647);
  nand g2126 (n_2504, n_1646, n_1648);
  nand g2127 (n_142, n_2502, n_2503, n_2504);
  xor g2128 (n_1656, n_1649, n_1650);
  and g2129 (n_1670, n_1649, n_1650);
  xor g2130 (n_2505, n_1651, n_1652);
  xor g2131 (n_1659, n_2505, n_1653);
  nand g2132 (n_2506, n_1651, n_1652);
  nand g2133 (n_2507, n_1653, n_1652);
  nand g2134 (n_2508, n_1651, n_1653);
  nand g2135 (n_1671, n_2506, n_2507, n_2508);
  xor g2136 (n_2509, n_1654, n_1655);
  xor g2137 (n_1660, n_2509, n_1656);
  nand g2138 (n_2510, n_1654, n_1655);
  nand g2139 (n_2511, n_1656, n_1655);
  nand g2140 (n_2512, n_1654, n_1656);
  nand g2141 (n_1673, n_2510, n_2511, n_2512);
  xor g2142 (n_2513, n_1657, n_1658);
  xor g2143 (n_1662, n_2513, n_1659);
  nand g2144 (n_2514, n_1657, n_1658);
  nand g2145 (n_2515, n_1659, n_1658);
  nand g2146 (n_2516, n_1657, n_1659);
  nand g2147 (n_1675, n_2514, n_2515, n_2516);
  xor g2148 (n_2517, n_1660, n_1661);
  xor g2149 (n_194, n_2517, n_1662);
  nand g2150 (n_2518, n_1660, n_1661);
  nand g2151 (n_2519, n_1662, n_1661);
  nand g2152 (n_2520, n_1660, n_1662);
  nand g2153 (n_141, n_2518, n_2519, n_2520);
  xor g2154 (n_1669, n_1663, n_1664);
  and g2155 (n_1685, n_1663, n_1664);
  xor g2156 (n_2521, n_1665, n_1666);
  xor g2157 (n_1672, n_2521, n_1667);
  nand g2158 (n_2522, n_1665, n_1666);
  nand g2159 (n_2523, n_1667, n_1666);
  nand g2160 (n_2524, n_1665, n_1667);
  nand g2161 (n_1687, n_2522, n_2523, n_2524);
  xor g2162 (n_2525, n_1668, n_1669);
  xor g2163 (n_1674, n_2525, n_1670);
  nand g2164 (n_2526, n_1668, n_1669);
  nand g2165 (n_2527, n_1670, n_1669);
  nand g2166 (n_2528, n_1668, n_1670);
  nand g2167 (n_1690, n_2526, n_2527, n_2528);
  xor g2168 (n_2529, n_1671, n_1672);
  xor g2169 (n_1676, n_2529, n_1673);
  nand g2170 (n_2530, n_1671, n_1672);
  nand g2171 (n_2531, n_1673, n_1672);
  nand g2172 (n_2532, n_1671, n_1673);
  nand g2173 (n_1693, n_2530, n_2531, n_2532);
  xor g2174 (n_2533, n_1674, n_1675);
  xor g2175 (n_193, n_2533, n_1676);
  nand g2176 (n_2534, n_1674, n_1675);
  nand g2177 (n_2535, n_1676, n_1675);
  nand g2178 (n_2536, n_1674, n_1676);
  nand g2179 (n_140, n_2534, n_2535, n_2536);
  xor g2180 (n_1686, n_1677, n_1678);
  and g2181 (n_1702, n_1677, n_1678);
  xor g2182 (n_2537, n_1679, n_1680);
  xor g2183 (n_1689, n_2537, n_1681);
  nand g2184 (n_2538, n_1679, n_1680);
  nand g2185 (n_2539, n_1681, n_1680);
  nand g2186 (n_2540, n_1679, n_1681);
  nand g2187 (n_1703, n_2538, n_2539, n_2540);
  xor g2188 (n_2541, n_1682, n_1683);
  xor g2189 (n_1688, n_2541, n_1684);
  nand g2190 (n_2542, n_1682, n_1683);
  nand g2191 (n_2543, n_1684, n_1683);
  nand g2192 (n_2544, n_1682, n_1684);
  nand g2193 (n_1704, n_2542, n_2543, n_2544);
  xor g2194 (n_2545, n_1685, n_1686);
  xor g2195 (n_1691, n_2545, n_1687);
  nand g2196 (n_2546, n_1685, n_1686);
  nand g2197 (n_2547, n_1687, n_1686);
  nand g2198 (n_2548, n_1685, n_1687);
  nand g2199 (n_1707, n_2546, n_2547, n_2548);
  xor g2200 (n_2549, n_1688, n_1689);
  xor g2201 (n_1692, n_2549, n_1690);
  nand g2202 (n_2550, n_1688, n_1689);
  nand g2203 (n_2551, n_1690, n_1689);
  nand g2204 (n_2552, n_1688, n_1690);
  nand g2205 (n_1709, n_2550, n_2551, n_2552);
  xor g2206 (n_2553, n_1691, n_1692);
  xor g2207 (n_192, n_2553, n_1693);
  nand g2208 (n_2554, n_1691, n_1692);
  nand g2209 (n_2555, n_1693, n_1692);
  nand g2210 (n_2556, n_1691, n_1693);
  nand g2211 (n_139, n_2554, n_2555, n_2556);
  xor g2212 (n_1701, n_1694, n_1695);
  and g2213 (n_1721, n_1694, n_1695);
  xor g2214 (n_2557, n_1696, n_1697);
  xor g2215 (n_1705, n_2557, n_1698);
  nand g2216 (n_2558, n_1696, n_1697);
  nand g2217 (n_2559, n_1698, n_1697);
  nand g2218 (n_2560, n_1696, n_1698);
  nand g2219 (n_1722, n_2558, n_2559, n_2560);
  xor g2220 (n_2561, n_1699, n_1700);
  xor g2221 (n_1706, n_2561, n_1701);
  nand g2222 (n_2562, n_1699, n_1700);
  nand g2223 (n_2563, n_1701, n_1700);
  nand g2224 (n_2564, n_1699, n_1701);
  nand g2225 (n_1725, n_2562, n_2563, n_2564);
  xor g2226 (n_2565, n_1702, n_1703);
  xor g2227 (n_1708, n_2565, n_1704);
  nand g2228 (n_2566, n_1702, n_1703);
  nand g2229 (n_2567, n_1704, n_1703);
  nand g2230 (n_2568, n_1702, n_1704);
  nand g2231 (n_1727, n_2566, n_2567, n_2568);
  xor g2232 (n_2569, n_1705, n_1706);
  xor g2233 (n_1710, n_2569, n_1707);
  nand g2234 (n_2570, n_1705, n_1706);
  nand g2235 (n_2571, n_1707, n_1706);
  nand g2236 (n_2572, n_1705, n_1707);
  nand g2237 (n_1729, n_2570, n_2571, n_2572);
  xor g2238 (n_2573, n_1708, n_1709);
  xor g2239 (n_191, n_2573, n_1710);
  nand g2240 (n_2574, n_1708, n_1709);
  nand g2241 (n_2575, n_1710, n_1709);
  nand g2242 (n_2576, n_1708, n_1710);
  nand g2243 (n_138, n_2574, n_2575, n_2576);
  xor g2244 (n_1720, n_1711, n_1712);
  and g2245 (n_1739, n_1711, n_1712);
  xor g2246 (n_2577, n_1713, n_1714);
  xor g2247 (n_1724, n_2577, n_1715);
  nand g2248 (n_2578, n_1713, n_1714);
  nand g2249 (n_2579, n_1715, n_1714);
  nand g2250 (n_2580, n_1713, n_1715);
  nand g2251 (n_1741, n_2578, n_2579, n_2580);
  xor g2252 (n_2581, n_1716, n_1717);
  xor g2253 (n_1723, n_2581, n_1718);
  nand g2254 (n_2582, n_1716, n_1717);
  nand g2255 (n_2583, n_1718, n_1717);
  nand g2256 (n_2584, n_1716, n_1718);
  nand g2257 (n_1742, n_2582, n_2583, n_2584);
  xor g2258 (n_2585, n_1719, n_1720);
  xor g2259 (n_1726, n_2585, n_1721);
  nand g2260 (n_2586, n_1719, n_1720);
  nand g2261 (n_2587, n_1721, n_1720);
  nand g2262 (n_2588, n_1719, n_1721);
  nand g2263 (n_1745, n_2586, n_2587, n_2588);
  xor g2264 (n_2589, n_1722, n_1723);
  xor g2265 (n_1728, n_2589, n_1724);
  nand g2266 (n_2590, n_1722, n_1723);
  nand g2267 (n_2591, n_1724, n_1723);
  nand g2268 (n_2592, n_1722, n_1724);
  nand g2269 (n_1747, n_2590, n_2591, n_2592);
  xor g2270 (n_2593, n_1725, n_1726);
  xor g2271 (n_1730, n_2593, n_1727);
  nand g2272 (n_2594, n_1725, n_1726);
  nand g2273 (n_2595, n_1727, n_1726);
  nand g2274 (n_2596, n_1725, n_1727);
  nand g2275 (n_1749, n_2594, n_2595, n_2596);
  xor g2276 (n_2597, n_1728, n_1729);
  xor g2277 (n_190, n_2597, n_1730);
  nand g2278 (n_2598, n_1728, n_1729);
  nand g2279 (n_2599, n_1730, n_1729);
  nand g2280 (n_2600, n_1728, n_1730);
  nand g2281 (n_137, n_2598, n_2599, n_2600);
  xor g2282 (n_1740, n_1731, n_1732);
  and g2283 (n_1762, n_1731, n_1732);
  xor g2284 (n_2601, n_1733, n_1734);
  xor g2285 (n_1744, n_2601, n_1735);
  nand g2286 (n_2602, n_1733, n_1734);
  nand g2287 (n_2603, n_1735, n_1734);
  nand g2288 (n_2604, n_1733, n_1735);
  nand g2289 (n_1763, n_2602, n_2603, n_2604);
  xor g2290 (n_2605, n_1736, n_1737);
  xor g2291 (n_1743, n_2605, n_1738);
  nand g2292 (n_2606, n_1736, n_1737);
  nand g2293 (n_2607, n_1738, n_1737);
  nand g2294 (n_2608, n_1736, n_1738);
  nand g2295 (n_1764, n_2606, n_2607, n_2608);
  xor g2296 (n_2609, n_1739, n_1740);
  xor g2297 (n_1746, n_2609, n_1741);
  nand g2298 (n_2610, n_1739, n_1740);
  nand g2299 (n_2611, n_1741, n_1740);
  nand g2300 (n_2612, n_1739, n_1741);
  nand g2301 (n_1768, n_2610, n_2611, n_2612);
  xor g2302 (n_2613, n_1742, n_1743);
  xor g2303 (n_1748, n_2613, n_1744);
  nand g2304 (n_2614, n_1742, n_1743);
  nand g2305 (n_2615, n_1744, n_1743);
  nand g2306 (n_2616, n_1742, n_1744);
  nand g2307 (n_1770, n_2614, n_2615, n_2616);
  xor g2308 (n_2617, n_1745, n_1746);
  xor g2309 (n_1750, n_2617, n_1747);
  nand g2310 (n_2618, n_1745, n_1746);
  nand g2311 (n_2619, n_1747, n_1746);
  nand g2312 (n_2620, n_1745, n_1747);
  nand g2313 (n_1772, n_2618, n_2619, n_2620);
  xor g2314 (n_2621, n_1748, n_1749);
  xor g2315 (n_189, n_2621, n_1750);
  nand g2316 (n_2622, n_1748, n_1749);
  nand g2317 (n_2623, n_1750, n_1749);
  nand g2318 (n_2624, n_1748, n_1750);
  nand g2319 (n_136, n_2622, n_2623, n_2624);
  xor g2320 (n_1761, n_1751, n_1752);
  and g2321 (n_1784, n_1751, n_1752);
  xor g2322 (n_2625, n_1753, n_1754);
  xor g2323 (n_1765, n_2625, n_1755);
  nand g2324 (n_2626, n_1753, n_1754);
  nand g2325 (n_2627, n_1755, n_1754);
  nand g2326 (n_2628, n_1753, n_1755);
  nand g2327 (n_1785, n_2626, n_2627, n_2628);
  xor g2328 (n_2629, n_1756, n_1757);
  xor g2329 (n_1766, n_2629, n_1758);
  nand g2330 (n_2630, n_1756, n_1757);
  nand g2331 (n_2631, n_1758, n_1757);
  nand g2332 (n_2632, n_1756, n_1758);
  nand g2333 (n_1786, n_2630, n_2631, n_2632);
  xor g2334 (n_2633, n_1759, n_1760);
  xor g2335 (n_1767, n_2633, n_1761);
  nand g2336 (n_2634, n_1759, n_1760);
  nand g2337 (n_2635, n_1761, n_1760);
  nand g2338 (n_2636, n_1759, n_1761);
  nand g2339 (n_1789, n_2634, n_2635, n_2636);
  xor g2340 (n_2637, n_1762, n_1763);
  xor g2341 (n_1769, n_2637, n_1764);
  nand g2342 (n_2638, n_1762, n_1763);
  nand g2343 (n_2639, n_1764, n_1763);
  nand g2344 (n_2640, n_1762, n_1764);
  nand g2345 (n_1790, n_2638, n_2639, n_2640);
  xor g2346 (n_2641, n_1765, n_1766);
  xor g2347 (n_1771, n_2641, n_1767);
  nand g2348 (n_2642, n_1765, n_1766);
  nand g2349 (n_2643, n_1767, n_1766);
  nand g2350 (n_2644, n_1765, n_1767);
  nand g2351 (n_1793, n_2642, n_2643, n_2644);
  xor g2352 (n_2645, n_1768, n_1769);
  xor g2353 (n_1773, n_2645, n_1770);
  nand g2354 (n_2646, n_1768, n_1769);
  nand g2355 (n_2647, n_1770, n_1769);
  nand g2356 (n_2648, n_1768, n_1770);
  nand g2357 (n_1795, n_2646, n_2647, n_2648);
  xor g2358 (n_2649, n_1771, n_1772);
  xor g2359 (n_188, n_2649, n_1773);
  nand g2360 (n_2650, n_1771, n_1772);
  nand g2361 (n_2651, n_1773, n_1772);
  nand g2362 (n_2652, n_1771, n_1773);
  nand g2363 (n_135, n_2650, n_2651, n_2652);
  xor g2364 (n_1783, n_1774, n_1775);
  and g2365 (n_1809, n_1774, n_1775);
  xor g2366 (n_2653, n_1776, n_1777);
  xor g2367 (n_1788, n_2653, n_1778);
  nand g2368 (n_2654, n_1776, n_1777);
  nand g2369 (n_2655, n_1778, n_1777);
  nand g2370 (n_2656, n_1776, n_1778);
  nand g2371 (n_1811, n_2654, n_2655, n_2656);
  xor g2372 (n_2657, n_1779, n_1780);
  xor g2373 (n_1787, n_2657, n_1781);
  nand g2374 (n_2658, n_1779, n_1780);
  nand g2375 (n_2659, n_1781, n_1780);
  nand g2376 (n_2660, n_1779, n_1781);
  nand g2377 (n_1810, n_2658, n_2659, n_2660);
  xor g2378 (n_2661, n_1782, n_1783);
  xor g2379 (n_1791, n_2661, n_1784);
  nand g2380 (n_2662, n_1782, n_1783);
  nand g2381 (n_2663, n_1784, n_1783);
  nand g2382 (n_2664, n_1782, n_1784);
  nand g2383 (n_1815, n_2662, n_2663, n_2664);
  xor g2384 (n_2665, n_1785, n_1786);
  xor g2385 (n_1792, n_2665, n_1787);
  nand g2386 (n_2666, n_1785, n_1786);
  nand g2387 (n_2667, n_1787, n_1786);
  nand g2388 (n_2668, n_1785, n_1787);
  nand g2389 (n_1817, n_2666, n_2667, n_2668);
  xor g2390 (n_2669, n_1788, n_1789);
  xor g2391 (n_1794, n_2669, n_1790);
  nand g2392 (n_2670, n_1788, n_1789);
  nand g2393 (n_2671, n_1790, n_1789);
  nand g2394 (n_2672, n_1788, n_1790);
  nand g2395 (n_1820, n_2670, n_2671, n_2672);
  xor g2396 (n_2673, n_1791, n_1792);
  xor g2397 (n_1796, n_2673, n_1793);
  nand g2398 (n_2674, n_1791, n_1792);
  nand g2399 (n_2675, n_1793, n_1792);
  nand g2400 (n_2676, n_1791, n_1793);
  nand g2401 (n_1821, n_2674, n_2675, n_2676);
  xor g2402 (n_2677, n_1794, n_1795);
  xor g2403 (n_187, n_2677, n_1796);
  nand g2404 (n_2678, n_1794, n_1795);
  nand g2405 (n_2679, n_1796, n_1795);
  nand g2406 (n_2680, n_1794, n_1796);
  nand g2407 (n_134, n_2678, n_2679, n_2680);
  xor g2408 (n_1808, n_1797, n_1798);
  and g2409 (n_1834, n_1797, n_1798);
  xor g2410 (n_2681, n_1799, n_1800);
  xor g2411 (n_1813, n_2681, n_1801);
  nand g2412 (n_2682, n_1799, n_1800);
  nand g2413 (n_2683, n_1801, n_1800);
  nand g2414 (n_2684, n_1799, n_1801);
  nand g2415 (n_1837, n_2682, n_2683, n_2684);
  xor g2416 (n_2685, n_1802, n_1803);
  xor g2417 (n_1814, n_2685, n_1804);
  nand g2418 (n_2686, n_1802, n_1803);
  nand g2419 (n_2687, n_1804, n_1803);
  nand g2420 (n_2688, n_1802, n_1804);
  nand g2421 (n_1835, n_2686, n_2687, n_2688);
  xor g2422 (n_2689, n_1805, n_1806);
  xor g2423 (n_1812, n_2689, n_1807);
  nand g2424 (n_2690, n_1805, n_1806);
  nand g2425 (n_2691, n_1807, n_1806);
  nand g2426 (n_2692, n_1805, n_1807);
  nand g2427 (n_1836, n_2690, n_2691, n_2692);
  xor g2428 (n_2693, n_1808, n_1809);
  xor g2429 (n_1816, n_2693, n_1810);
  nand g2430 (n_2694, n_1808, n_1809);
  nand g2431 (n_2695, n_1810, n_1809);
  nand g2432 (n_2696, n_1808, n_1810);
  nand g2433 (n_1841, n_2694, n_2695, n_2696);
  xor g2434 (n_2697, n_1811, n_1812);
  xor g2435 (n_1818, n_2697, n_1813);
  nand g2436 (n_2698, n_1811, n_1812);
  nand g2437 (n_2699, n_1813, n_1812);
  nand g2438 (n_2700, n_1811, n_1813);
  nand g2439 (n_1842, n_2698, n_2699, n_2700);
  xor g2440 (n_2701, n_1814, n_1815);
  xor g2441 (n_1819, n_2701, n_1816);
  nand g2442 (n_2702, n_1814, n_1815);
  nand g2443 (n_2703, n_1816, n_1815);
  nand g2444 (n_2704, n_1814, n_1816);
  nand g2445 (n_1845, n_2702, n_2703, n_2704);
  xor g2446 (n_2705, n_1817, n_1818);
  xor g2447 (n_1822, n_2705, n_1819);
  nand g2448 (n_2706, n_1817, n_1818);
  nand g2449 (n_2707, n_1819, n_1818);
  nand g2450 (n_2708, n_1817, n_1819);
  nand g2451 (n_1848, n_2706, n_2707, n_2708);
  xor g2452 (n_2709, n_1820, n_1821);
  xor g2453 (n_186, n_2709, n_1822);
  nand g2454 (n_2710, n_1820, n_1821);
  nand g2455 (n_2711, n_1822, n_1821);
  nand g2456 (n_2712, n_1820, n_1822);
  nand g2457 (n_133, n_2710, n_2711, n_2712);
  xor g2458 (n_1833, n_1823, n_1824);
  and g2459 (n_1862, n_1823, n_1824);
  xor g2460 (n_2713, n_1825, n_1826);
  xor g2461 (n_1838, n_2713, n_1827);
  nand g2462 (n_2714, n_1825, n_1826);
  nand g2463 (n_2715, n_1827, n_1826);
  nand g2464 (n_2716, n_1825, n_1827);
  nand g2465 (n_1864, n_2714, n_2715, n_2716);
  xor g2466 (n_2717, n_1828, n_1829);
  xor g2467 (n_1839, n_2717, n_1830);
  nand g2468 (n_2718, n_1828, n_1829);
  nand g2469 (n_2719, n_1830, n_1829);
  nand g2470 (n_2720, n_1828, n_1830);
  nand g2471 (n_1863, n_2718, n_2719, n_2720);
  xor g2472 (n_2721, n_1831, n_1832);
  xor g2473 (n_1840, n_2721, n_1833);
  nand g2474 (n_2722, n_1831, n_1832);
  nand g2475 (n_2723, n_1833, n_1832);
  nand g2476 (n_2724, n_1831, n_1833);
  nand g2477 (n_1868, n_2722, n_2723, n_2724);
  xor g2478 (n_2725, n_1834, n_1835);
  xor g2479 (n_1843, n_2725, n_1836);
  nand g2480 (n_2726, n_1834, n_1835);
  nand g2481 (n_2727, n_1836, n_1835);
  nand g2482 (n_2728, n_1834, n_1836);
  nand g2483 (n_1870, n_2726, n_2727, n_2728);
  xor g2484 (n_2729, n_1837, n_1838);
  xor g2485 (n_1844, n_2729, n_1839);
  nand g2486 (n_2730, n_1837, n_1838);
  nand g2487 (n_2731, n_1839, n_1838);
  nand g2488 (n_2732, n_1837, n_1839);
  nand g2489 (n_1872, n_2730, n_2731, n_2732);
  xor g2490 (n_2733, n_1840, n_1841);
  xor g2491 (n_1846, n_2733, n_1842);
  nand g2492 (n_2734, n_1840, n_1841);
  nand g2493 (n_2735, n_1842, n_1841);
  nand g2494 (n_2736, n_1840, n_1842);
  nand g2495 (n_1875, n_2734, n_2735, n_2736);
  xor g2496 (n_2737, n_1843, n_1844);
  xor g2497 (n_1847, n_2737, n_1845);
  nand g2498 (n_2738, n_1843, n_1844);
  nand g2499 (n_2739, n_1845, n_1844);
  nand g2500 (n_2740, n_1843, n_1845);
  nand g2501 (n_1876, n_2738, n_2739, n_2740);
  xor g2502 (n_2741, n_1846, n_1847);
  xor g2503 (n_185, n_2741, n_1848);
  nand g2504 (n_2742, n_1846, n_1847);
  nand g2505 (n_2743, n_1848, n_1847);
  nand g2506 (n_2744, n_1846, n_1848);
  nand g2507 (n_132, n_2742, n_2743, n_2744);
  xor g2508 (n_1861, n_1849, n_1850);
  and g2509 (n_1890, n_1849, n_1850);
  xor g2510 (n_2745, n_1851, n_1852);
  xor g2511 (n_1866, n_2745, n_1853);
  nand g2512 (n_2746, n_1851, n_1852);
  nand g2513 (n_2747, n_1853, n_1852);
  nand g2514 (n_2748, n_1851, n_1853);
  nand g2515 (n_1892, n_2746, n_2747, n_2748);
  xor g2516 (n_2749, n_1854, n_1855);
  xor g2517 (n_1867, n_2749, n_1856);
  nand g2518 (n_2750, n_1854, n_1855);
  nand g2519 (n_2751, n_1856, n_1855);
  nand g2520 (n_2752, n_1854, n_1856);
  nand g2521 (n_1893, n_2750, n_2751, n_2752);
  xor g2522 (n_2753, n_1857, n_1858);
  xor g2523 (n_1865, n_2753, n_1859);
  nand g2524 (n_2754, n_1857, n_1858);
  nand g2525 (n_2755, n_1859, n_1858);
  nand g2526 (n_2756, n_1857, n_1859);
  nand g2527 (n_1891, n_2754, n_2755, n_2756);
  xor g2528 (n_2757, n_1860, n_1861);
  xor g2529 (n_1869, n_2757, n_1862);
  nand g2530 (n_2758, n_1860, n_1861);
  nand g2531 (n_2759, n_1862, n_1861);
  nand g2532 (n_2760, n_1860, n_1862);
  nand g2533 (n_1897, n_2758, n_2759, n_2760);
  xor g2534 (n_2761, n_1863, n_1864);
  xor g2535 (n_1871, n_2761, n_1865);
  nand g2536 (n_2762, n_1863, n_1864);
  nand g2537 (n_2763, n_1865, n_1864);
  nand g2538 (n_2764, n_1863, n_1865);
  nand g2539 (n_1899, n_2762, n_2763, n_2764);
  xor g2540 (n_2765, n_1866, n_1867);
  xor g2541 (n_1873, n_2765, n_1868);
  nand g2542 (n_2766, n_1866, n_1867);
  nand g2543 (n_2767, n_1868, n_1867);
  nand g2544 (n_2768, n_1866, n_1868);
  nand g2545 (n_1902, n_2766, n_2767, n_2768);
  xor g2546 (n_2769, n_1869, n_1870);
  xor g2547 (n_1874, n_2769, n_1871);
  nand g2548 (n_2770, n_1869, n_1870);
  nand g2549 (n_2771, n_1871, n_1870);
  nand g2550 (n_2772, n_1869, n_1871);
  nand g2551 (n_1903, n_2770, n_2771, n_2772);
  xor g2552 (n_2773, n_1872, n_1873);
  xor g2553 (n_1877, n_2773, n_1874);
  nand g2554 (n_2774, n_1872, n_1873);
  nand g2555 (n_2775, n_1874, n_1873);
  nand g2556 (n_2776, n_1872, n_1874);
  nand g2557 (n_1906, n_2774, n_2775, n_2776);
  xor g2558 (n_2777, n_1875, n_1876);
  xor g2559 (n_184, n_2777, n_1877);
  nand g2560 (n_2778, n_1875, n_1876);
  nand g2561 (n_2779, n_1877, n_1876);
  nand g2562 (n_2780, n_1875, n_1877);
  nand g2563 (n_131, n_2778, n_2779, n_2780);
  xor g2564 (n_1889, n_1878, n_1879);
  and g2565 (n_1921, n_1878, n_1879);
  xor g2566 (n_2781, n_1880, n_1881);
  xor g2567 (n_1894, n_2781, n_1882);
  nand g2568 (n_2782, n_1880, n_1881);
  nand g2569 (n_2783, n_1882, n_1881);
  nand g2570 (n_2784, n_1880, n_1882);
  nand g2571 (n_1924, n_2782, n_2783, n_2784);
  xor g2572 (n_2785, n_1883, n_1884);
  xor g2573 (n_1895, n_2785, n_1885);
  nand g2574 (n_2786, n_1883, n_1884);
  nand g2575 (n_2787, n_1885, n_1884);
  nand g2576 (n_2788, n_1883, n_1885);
  nand g2577 (n_1922, n_2786, n_2787, n_2788);
  xor g2578 (n_2789, n_1886, n_1887);
  xor g2579 (n_1896, n_2789, n_1888);
  nand g2580 (n_2790, n_1886, n_1887);
  nand g2581 (n_2791, n_1888, n_1887);
  nand g2582 (n_2792, n_1886, n_1888);
  nand g2583 (n_1923, n_2790, n_2791, n_2792);
  xor g2584 (n_2793, n_1889, n_1890);
  xor g2585 (n_1898, n_2793, n_1891);
  nand g2586 (n_2794, n_1889, n_1890);
  nand g2587 (n_2795, n_1891, n_1890);
  nand g2588 (n_2796, n_1889, n_1891);
  nand g2589 (n_1929, n_2794, n_2795, n_2796);
  xor g2590 (n_2797, n_1892, n_1893);
  xor g2591 (n_1900, n_2797, n_1894);
  nand g2592 (n_2798, n_1892, n_1893);
  nand g2593 (n_2799, n_1894, n_1893);
  nand g2594 (n_2800, n_1892, n_1894);
  nand g2595 (n_1931, n_2798, n_2799, n_2800);
  xor g2596 (n_2801, n_1895, n_1896);
  xor g2597 (n_1901, n_2801, n_1897);
  nand g2598 (n_2802, n_1895, n_1896);
  nand g2599 (n_2803, n_1897, n_1896);
  nand g2600 (n_2804, n_1895, n_1897);
  nand g2601 (n_1932, n_2802, n_2803, n_2804);
  xor g2602 (n_2805, n_1898, n_1899);
  xor g2603 (n_1904, n_2805, n_1900);
  nand g2604 (n_2806, n_1898, n_1899);
  nand g2605 (n_2807, n_1900, n_1899);
  nand g2606 (n_2808, n_1898, n_1900);
  nand g2607 (n_1935, n_2806, n_2807, n_2808);
  xor g2608 (n_2809, n_1901, n_1902);
  xor g2609 (n_1905, n_2809, n_1903);
  nand g2610 (n_2810, n_1901, n_1902);
  nand g2611 (n_2811, n_1903, n_1902);
  nand g2612 (n_2812, n_1901, n_1903);
  nand g2613 (n_1938, n_2810, n_2811, n_2812);
  xor g2614 (n_2813, n_1904, n_1905);
  xor g2615 (n_183, n_2813, n_1906);
  nand g2616 (n_2814, n_1904, n_1905);
  nand g2617 (n_2815, n_1906, n_1905);
  nand g2618 (n_2816, n_1904, n_1906);
  nand g2619 (n_130, n_2814, n_2815, n_2816);
  xor g2620 (n_1920, n_1907, n_1908);
  and g2621 (n_1952, n_1907, n_1908);
  xor g2622 (n_2817, n_1909, n_1910);
  xor g2623 (n_1927, n_2817, n_1911);
  nand g2624 (n_2818, n_1909, n_1910);
  nand g2625 (n_2819, n_1911, n_1910);
  nand g2626 (n_2820, n_1909, n_1911);
  nand g2627 (n_1954, n_2818, n_2819, n_2820);
  xor g2628 (n_2821, n_1912, n_1913);
  xor g2629 (n_1926, n_2821, n_1914);
  nand g2630 (n_2822, n_1912, n_1913);
  nand g2631 (n_2823, n_1914, n_1913);
  nand g2632 (n_2824, n_1912, n_1914);
  nand g2633 (n_1955, n_2822, n_2823, n_2824);
  xor g2634 (n_2825, n_1915, n_1916);
  xor g2635 (n_1925, n_2825, n_1917);
  nand g2636 (n_2826, n_1915, n_1916);
  nand g2637 (n_2827, n_1917, n_1916);
  nand g2638 (n_2828, n_1915, n_1917);
  nand g2639 (n_1953, n_2826, n_2827, n_2828);
  xor g2640 (n_2829, n_1918, n_1919);
  xor g2641 (n_1928, n_2829, n_1920);
  nand g2642 (n_2830, n_1918, n_1919);
  nand g2643 (n_2831, n_1920, n_1919);
  nand g2644 (n_2832, n_1918, n_1920);
  nand g2645 (n_1959, n_2830, n_2831, n_2832);
  xor g2646 (n_2833, n_1921, n_1922);
  xor g2647 (n_1930, n_2833, n_1923);
  nand g2648 (n_2834, n_1921, n_1922);
  nand g2649 (n_2835, n_1923, n_1922);
  nand g2650 (n_2836, n_1921, n_1923);
  nand g2651 (n_1960, n_2834, n_2835, n_2836);
  xor g2652 (n_2837, n_1924, n_1925);
  xor g2653 (n_1933, n_2837, n_1926);
  nand g2654 (n_2838, n_1924, n_1925);
  nand g2655 (n_2839, n_1926, n_1925);
  nand g2656 (n_2840, n_1924, n_1926);
  nand g2657 (n_1962, n_2838, n_2839, n_2840);
  xor g2658 (n_2841, n_1927, n_1928);
  xor g2659 (n_1934, n_2841, n_1929);
  nand g2660 (n_2842, n_1927, n_1928);
  nand g2661 (n_2843, n_1929, n_1928);
  nand g2662 (n_2844, n_1927, n_1929);
  nand g2663 (n_1965, n_2842, n_2843, n_2844);
  xor g2664 (n_2845, n_1930, n_1931);
  xor g2665 (n_1936, n_2845, n_1932);
  nand g2666 (n_2846, n_1930, n_1931);
  nand g2667 (n_2847, n_1932, n_1931);
  nand g2668 (n_2848, n_1930, n_1932);
  nand g2669 (n_1967, n_2846, n_2847, n_2848);
  xor g2670 (n_2849, n_1933, n_1934);
  xor g2671 (n_1937, n_2849, n_1935);
  nand g2672 (n_2850, n_1933, n_1934);
  nand g2673 (n_2851, n_1935, n_1934);
  nand g2674 (n_2852, n_1933, n_1935);
  nand g2675 (n_1969, n_2850, n_2851, n_2852);
  xor g2676 (n_2853, n_1936, n_1937);
  xor g2677 (n_182, n_2853, n_1938);
  nand g2678 (n_2854, n_1936, n_1937);
  nand g2679 (n_2855, n_1938, n_1937);
  nand g2680 (n_2856, n_1936, n_1938);
  nand g2681 (n_129, n_2854, n_2855, n_2856);
  xor g2682 (n_1951, n_1939, n_1940);
  and g2683 (n_1984, n_1939, n_1940);
  xor g2684 (n_2857, n_1941, n_1942);
  xor g2685 (n_1958, n_2857, n_1943);
  nand g2686 (n_2858, n_1941, n_1942);
  nand g2687 (n_2859, n_1943, n_1942);
  nand g2688 (n_2860, n_1941, n_1943);
  nand g2689 (n_1987, n_2858, n_2859, n_2860);
  xor g2690 (n_2861, n_1944, n_1945);
  xor g2691 (n_1957, n_2861, n_1946);
  nand g2692 (n_2862, n_1944, n_1945);
  nand g2693 (n_2863, n_1946, n_1945);
  nand g2694 (n_2864, n_1944, n_1946);
  nand g2695 (n_1985, n_2862, n_2863, n_2864);
  xor g2696 (n_2865, n_1947, n_1948);
  xor g2697 (n_1956, n_2865, n_1949);
  nand g2698 (n_2866, n_1947, n_1948);
  nand g2699 (n_2867, n_1949, n_1948);
  nand g2700 (n_2868, n_1947, n_1949);
  nand g2701 (n_1986, n_2866, n_2867, n_2868);
  xor g2702 (n_2869, n_1950, n_1951);
  xor g2703 (n_1961, n_2869, n_1952);
  nand g2704 (n_2870, n_1950, n_1951);
  nand g2705 (n_2871, n_1952, n_1951);
  nand g2706 (n_2872, n_1950, n_1952);
  nand g2707 (n_1992, n_2870, n_2871, n_2872);
  xor g2708 (n_2873, n_1953, n_1954);
  xor g2709 (n_1963, n_2873, n_1955);
  nand g2710 (n_2874, n_1953, n_1954);
  nand g2711 (n_2875, n_1955, n_1954);
  nand g2712 (n_2876, n_1953, n_1955);
  nand g2713 (n_1993, n_2874, n_2875, n_2876);
  xor g2714 (n_2877, n_1956, n_1957);
  xor g2715 (n_1964, n_2877, n_1958);
  nand g2716 (n_2878, n_1956, n_1957);
  nand g2717 (n_2879, n_1958, n_1957);
  nand g2718 (n_2880, n_1956, n_1958);
  nand g2719 (n_1996, n_2878, n_2879, n_2880);
  xor g2720 (n_2881, n_1959, n_1960);
  xor g2721 (n_1966, n_2881, n_1961);
  nand g2722 (n_2882, n_1959, n_1960);
  nand g2723 (n_2883, n_1961, n_1960);
  nand g2724 (n_2884, n_1959, n_1961);
  nand g2725 (n_1998, n_2882, n_2883, n_2884);
  xor g2726 (n_2885, n_1962, n_1963);
  xor g2727 (n_1968, n_2885, n_1964);
  nand g2728 (n_2886, n_1962, n_1963);
  nand g2729 (n_2887, n_1964, n_1963);
  nand g2730 (n_2888, n_1962, n_1964);
  nand g2731 (n_2000, n_2886, n_2887, n_2888);
  xor g2732 (n_2889, n_1965, n_1966);
  xor g2733 (n_1970, n_2889, n_1967);
  nand g2734 (n_2890, n_1965, n_1966);
  nand g2735 (n_2891, n_1967, n_1966);
  nand g2736 (n_2892, n_1965, n_1967);
  nand g2737 (n_2003, n_2890, n_2891, n_2892);
  xor g2738 (n_2893, n_1968, n_1969);
  xor g2739 (n_181, n_2893, n_1970);
  nand g2740 (n_2894, n_1968, n_1969);
  nand g2741 (n_2895, n_1970, n_1969);
  nand g2742 (n_2896, n_1968, n_1970);
  nand g2743 (n_128, n_2894, n_2895, n_2896);
  xor g2745 (n_1990, n_2897, n_1973);
  nand g2747 (n_2899, n_1973, n_1972);
  nand g2749 (n_2020, n_2898, n_2899, n_2900);
  xor g2750 (n_2901, n_1974, n_1975);
  xor g2751 (n_1991, n_2901, n_1976);
  nand g2752 (n_2902, n_1974, n_1975);
  nand g2753 (n_2903, n_1976, n_1975);
  nand g2754 (n_2904, n_1974, n_1976);
  nand g2755 (n_2019, n_2902, n_2903, n_2904);
  xor g2756 (n_2905, n_1977, n_1978);
  xor g2757 (n_1989, n_2905, n_1979);
  nand g2758 (n_2906, n_1977, n_1978);
  nand g2759 (n_2907, n_1979, n_1978);
  nand g2760 (n_2908, n_1977, n_1979);
  nand g2761 (n_2021, n_2906, n_2907, n_2908);
  xor g2762 (n_2909, n_1980, n_1981);
  xor g2763 (n_1988, n_2909, n_1982);
  nand g2764 (n_2910, n_1980, n_1981);
  nand g2765 (n_2911, n_1982, n_1981);
  nand g2766 (n_2912, n_1980, n_1982);
  nand g2767 (n_2022, n_2910, n_2911, n_2912);
  xor g2768 (n_2913, n_1983, n_1984);
  xor g2769 (n_1994, n_2913, n_1985);
  nand g2770 (n_2914, n_1983, n_1984);
  nand g2771 (n_2915, n_1985, n_1984);
  nand g2772 (n_2916, n_1983, n_1985);
  nand g2773 (n_2027, n_2914, n_2915, n_2916);
  xor g2774 (n_2917, n_1986, n_1987);
  xor g2775 (n_1995, n_2917, n_1988);
  nand g2776 (n_2918, n_1986, n_1987);
  nand g2777 (n_2919, n_1988, n_1987);
  nand g2778 (n_2920, n_1986, n_1988);
  nand g2779 (n_2028, n_2918, n_2919, n_2920);
  xor g2780 (n_2921, n_1989, n_1990);
  xor g2781 (n_1997, n_2921, n_1991);
  nand g2782 (n_2922, n_1989, n_1990);
  nand g2783 (n_2923, n_1991, n_1990);
  nand g2784 (n_2924, n_1989, n_1991);
  nand g2785 (n_2030, n_2922, n_2923, n_2924);
  xor g2786 (n_2925, n_1992, n_1993);
  xor g2787 (n_1999, n_2925, n_1994);
  nand g2788 (n_2926, n_1992, n_1993);
  nand g2789 (n_2927, n_1994, n_1993);
  nand g2790 (n_2928, n_1992, n_1994);
  nand g2791 (n_2033, n_2926, n_2927, n_2928);
  xor g2792 (n_2929, n_1995, n_1996);
  xor g2793 (n_2001, n_2929, n_1997);
  nand g2794 (n_2930, n_1995, n_1996);
  nand g2795 (n_2931, n_1997, n_1996);
  nand g2796 (n_2932, n_1995, n_1997);
  nand g2797 (n_2035, n_2930, n_2931, n_2932);
  xor g2798 (n_2933, n_1998, n_1999);
  xor g2799 (n_2002, n_2933, n_2000);
  nand g2800 (n_2934, n_1998, n_1999);
  nand g2801 (n_2935, n_2000, n_1999);
  nand g2802 (n_2936, n_1998, n_2000);
  nand g2803 (n_2037, n_2934, n_2935, n_2936);
  xor g2804 (n_2937, n_2001, n_2002);
  xor g2805 (n_180, n_2937, n_2003);
  nand g2806 (n_2938, n_2001, n_2002);
  nand g2807 (n_2939, n_2003, n_2002);
  nand g2808 (n_2940, n_2001, n_2003);
  nand g2809 (n_127, n_2938, n_2939, n_2940);
  xor g2812 (n_2941, n_2006, n_2007);
  xor g2813 (n_2025, n_2941, n_2008);
  nand g2814 (n_2942, n_2006, n_2007);
  nand g2815 (n_2943, n_2008, n_2007);
  nand g2816 (n_2944, n_2006, n_2008);
  nand g2817 (n_2055, n_2942, n_2943, n_2944);
  xor g2818 (n_2945, n_2009, n_2010);
  xor g2819 (n_2026, n_2945, n_2011);
  nand g2820 (n_2946, n_2009, n_2010);
  nand g2821 (n_2947, n_2011, n_2010);
  nand g2822 (n_2948, n_2009, n_2011);
  nand g2823 (n_2056, n_2946, n_2947, n_2948);
  xor g2825 (n_2024, n_2949, n_2014);
  nand g2827 (n_2951, n_2014, n_2013);
  nand g2829 (n_2057, n_2950, n_2951, n_2952);
  xor g2830 (n_2953, n_2015, n_2016);
  xor g2831 (n_2023, n_2953, n_2017);
  nand g2832 (n_2954, n_2015, n_2016);
  nand g2833 (n_2955, n_2017, n_2016);
  nand g2834 (n_2956, n_2015, n_2017);
  nand g2835 (n_2054, n_2954, n_2955, n_2956);
  xor g2836 (n_2957, n_1501, n_2019);
  xor g2837 (n_2031, n_2957, n_2020);
  nand g2838 (n_2958, n_1501, n_2019);
  nand g2839 (n_2959, n_2020, n_2019);
  nand g2840 (n_2960, n_1501, n_2020);
  nand g2841 (n_2062, n_2958, n_2959, n_2960);
  xor g2842 (n_2961, n_2021, n_2022);
  xor g2843 (n_2029, n_2961, n_2023);
  nand g2844 (n_2962, n_2021, n_2022);
  nand g2845 (n_2963, n_2023, n_2022);
  nand g2846 (n_2964, n_2021, n_2023);
  nand g2847 (n_2065, n_2962, n_2963, n_2964);
  xor g2848 (n_2965, n_2024, n_2025);
  xor g2849 (n_2032, n_2965, n_2026);
  nand g2850 (n_2966, n_2024, n_2025);
  nand g2851 (n_2967, n_2026, n_2025);
  nand g2852 (n_2968, n_2024, n_2026);
  nand g2853 (n_2063, n_2966, n_2967, n_2968);
  xor g2854 (n_2969, n_2027, n_2028);
  xor g2855 (n_2036, n_2969, n_2029);
  nand g2856 (n_2970, n_2027, n_2028);
  nand g2857 (n_2971, n_2029, n_2028);
  nand g2858 (n_2972, n_2027, n_2029);
  nand g2859 (n_2068, n_2970, n_2971, n_2972);
  xor g2860 (n_2973, n_2030, n_2031);
  xor g2861 (n_2034, n_2973, n_2032);
  nand g2862 (n_2974, n_2030, n_2031);
  nand g2863 (n_2975, n_2032, n_2031);
  nand g2864 (n_2976, n_2030, n_2032);
  nand g2865 (n_2070, n_2974, n_2975, n_2976);
  xor g2866 (n_2977, n_2033, n_2034);
  xor g2867 (n_2038, n_2977, n_2035);
  nand g2868 (n_2978, n_2033, n_2034);
  nand g2869 (n_2979, n_2035, n_2034);
  nand g2870 (n_2980, n_2033, n_2035);
  nand g2871 (n_2072, n_2978, n_2979, n_2980);
  xor g2872 (n_2981, n_2036, n_2037);
  xor g2873 (n_179, n_2981, n_2038);
  nand g2874 (n_2982, n_2036, n_2037);
  nand g2875 (n_2983, n_2038, n_2037);
  nand g2876 (n_2984, n_2036, n_2038);
  nand g2877 (n_126, n_2982, n_2983, n_2984);
  xor g2880 (n_2985, n_2041, n_2042);
  xor g2881 (n_2060, n_2985, n_2043);
  nand g2882 (n_2986, n_2041, n_2042);
  nand g2883 (n_2987, n_2043, n_2042);
  nand g2884 (n_2988, n_2041, n_2043);
  nand g2885 (n_2089, n_2986, n_2987, n_2988);
  xor g2886 (n_2989, n_2044, n_2045);
  xor g2887 (n_2061, n_2989, n_2046);
  nand g2888 (n_2990, n_2044, n_2045);
  nand g2889 (n_2991, n_2046, n_2045);
  nand g2890 (n_2992, n_2044, n_2046);
  nand g2891 (n_2087, n_2990, n_2991, n_2992);
  xor g2892 (n_2993, n_2047, n_2048);
  xor g2893 (n_2059, n_2993, n_2049);
  nand g2894 (n_2994, n_2047, n_2048);
  nand g2895 (n_2995, n_2049, n_2048);
  nand g2896 (n_2996, n_2047, n_2049);
  nand g2897 (n_2088, n_2994, n_2995, n_2996);
  xor g2898 (n_2997, n_2050, n_2051);
  xor g2899 (n_2058, n_2997, n_1505);
  nand g2900 (n_2998, n_2050, n_2051);
  nand g2901 (n_2999, n_1505, n_2051);
  nand g2902 (n_3000, n_2050, n_1505);
  nand g2903 (n_2090, n_2998, n_2999, n_3000);
  xor g2905 (n_2066, n_3001, n_2055);
  nand g2907 (n_3003, n_2055, n_2054);
  nand g2909 (n_2095, n_3002, n_3003, n_3004);
  xor g2910 (n_3005, n_2056, n_2057);
  xor g2911 (n_2064, n_3005, n_2058);
  nand g2912 (n_3006, n_2056, n_2057);
  nand g2913 (n_3007, n_2058, n_2057);
  nand g2914 (n_3008, n_2056, n_2058);
  nand g2915 (n_2097, n_3006, n_3007, n_3008);
  xor g2916 (n_3009, n_2059, n_2060);
  xor g2917 (n_2067, n_3009, n_2061);
  nand g2918 (n_3010, n_2059, n_2060);
  nand g2919 (n_3011, n_2061, n_2060);
  nand g2920 (n_3012, n_2059, n_2061);
  nand g2921 (n_2096, n_3010, n_3011, n_3012);
  xor g2922 (n_3013, n_2062, n_2063);
  xor g2923 (n_2071, n_3013, n_2064);
  nand g2924 (n_3014, n_2062, n_2063);
  nand g2925 (n_3015, n_2064, n_2063);
  nand g2926 (n_3016, n_2062, n_2064);
  nand g2927 (n_2101, n_3014, n_3015, n_3016);
  xor g2928 (n_3017, n_2065, n_2066);
  xor g2929 (n_2069, n_3017, n_2067);
  nand g2930 (n_3018, n_2065, n_2066);
  nand g2931 (n_3019, n_2067, n_2066);
  nand g2932 (n_3020, n_2065, n_2067);
  nand g2933 (n_2103, n_3018, n_3019, n_3020);
  xor g2934 (n_3021, n_2068, n_2069);
  xor g2935 (n_2073, n_3021, n_2070);
  nand g2936 (n_3022, n_2068, n_2069);
  nand g2937 (n_3023, n_2070, n_2069);
  nand g2938 (n_3024, n_2068, n_2070);
  nand g2939 (n_2105, n_3022, n_3023, n_3024);
  xor g2940 (n_3025, n_2071, n_2072);
  xor g2941 (n_178, n_3025, n_2073);
  nand g2942 (n_3026, n_2071, n_2072);
  nand g2943 (n_3027, n_2073, n_2072);
  nand g2944 (n_3028, n_2071, n_2073);
  nand g2945 (n_125, n_3026, n_3027, n_3028);
  xor g2947 (n_2093, n_3029, n_2076);
  nand g2949 (n_3031, n_2076, n_2075);
  nand g2951 (n_2122, n_3030, n_3031, n_3032);
  xor g2953 (n_2094, n_3033, n_2079);
  nand g2955 (n_3035, n_2079, n_2078);
  nand g2957 (n_2120, n_3034, n_3035, n_3036);
  xor g2958 (n_3037, n_2080, n_2081);
  xor g2959 (n_2092, n_3037, n_2082);
  nand g2960 (n_3038, n_2080, n_2081);
  nand g2961 (n_3039, n_2082, n_2081);
  nand g2962 (n_3040, n_2080, n_2082);
  nand g2963 (n_2123, n_3038, n_3039, n_3040);
  xor g2964 (n_3041, n_2083, n_2084);
  xor g2965 (n_2091, n_3041, n_2085);
  nand g2966 (n_3042, n_2083, n_2084);
  nand g2967 (n_3043, n_2085, n_2084);
  nand g2968 (n_3044, n_2083, n_2085);
  nand g2969 (n_2121, n_3042, n_3043, n_3044);
  xor g2971 (n_2098, n_3045, n_2088);
  nand g2973 (n_3047, n_2088, n_2087);
  nand g2975 (n_2127, n_3046, n_3047, n_3048);
  xor g2976 (n_3049, n_2089, n_2090);
  xor g2977 (n_2100, n_3049, n_2091);
  nand g2978 (n_3050, n_2089, n_2090);
  nand g2979 (n_3051, n_2091, n_2090);
  nand g2980 (n_3052, n_2089, n_2091);
  nand g2981 (n_2129, n_3050, n_3051, n_3052);
  xor g2982 (n_3053, n_2092, n_2093);
  xor g2983 (n_2099, n_3053, n_2094);
  nand g2984 (n_3054, n_2092, n_2093);
  nand g2985 (n_3055, n_2094, n_2093);
  nand g2986 (n_3056, n_2092, n_2094);
  nand g2987 (n_2131, n_3054, n_3055, n_3056);
  xor g2988 (n_3057, n_2095, n_2096);
  xor g2989 (n_2102, n_3057, n_2097);
  nand g2990 (n_3058, n_2095, n_2096);
  nand g2991 (n_3059, n_2097, n_2096);
  nand g2992 (n_3060, n_2095, n_2097);
  nand g2993 (n_2133, n_3058, n_3059, n_3060);
  xor g2994 (n_3061, n_2098, n_2099);
  xor g2995 (n_2104, n_3061, n_2100);
  nand g2996 (n_3062, n_2098, n_2099);
  nand g2997 (n_3063, n_2100, n_2099);
  nand g2998 (n_3064, n_2098, n_2100);
  nand g2999 (n_2136, n_3062, n_3063, n_3064);
  xor g3000 (n_3065, n_2101, n_2102);
  xor g3001 (n_2106, n_3065, n_2103);
  nand g3002 (n_3066, n_2101, n_2102);
  nand g3003 (n_3067, n_2103, n_2102);
  nand g3004 (n_3068, n_2101, n_2103);
  nand g3005 (n_2138, n_3066, n_3067, n_3068);
  xor g3006 (n_3069, n_2104, n_2105);
  xor g3007 (n_177, n_3069, n_2106);
  nand g3008 (n_3070, n_2104, n_2105);
  nand g3009 (n_3071, n_2106, n_2105);
  nand g3010 (n_3072, n_2104, n_2106);
  nand g3011 (n_124, n_3070, n_3071, n_3072);
  xor g3014 (n_3073, n_2109, n_2110);
  xor g3015 (n_2126, n_3073, n_2111);
  nand g3016 (n_3074, n_2109, n_2110);
  nand g3017 (n_3075, n_2111, n_2110);
  nand g3018 (n_3076, n_2109, n_2111);
  nand g3019 (n_2153, n_3074, n_3075, n_3076);
  xor g3020 (n_3077, n_2112, n_2113);
  xor g3021 (n_2124, n_3077, n_2114);
  nand g3022 (n_3078, n_2112, n_2113);
  nand g3023 (n_3079, n_2114, n_2113);
  nand g3024 (n_3080, n_2112, n_2114);
  nand g3025 (n_2151, n_3078, n_3079, n_3080);
  xor g3026 (n_3081, n_2115, n_2116);
  xor g3027 (n_2125, n_3081, n_2117);
  nand g3028 (n_3082, n_2115, n_2116);
  nand g3029 (n_3083, n_2117, n_2116);
  nand g3030 (n_3084, n_2115, n_2117);
  nand g3031 (n_2152, n_3082, n_3083, n_3084);
  xor g3032 (n_3085, n_2118, n_1513);
  xor g3033 (n_2128, n_3085, n_2120);
  nand g3034 (n_3086, n_2118, n_1513);
  nand g3035 (n_3087, n_2120, n_1513);
  nand g3036 (n_3088, n_2118, n_2120);
  nand g3037 (n_2159, n_3086, n_3087, n_3088);
  xor g3038 (n_3089, n_2121, n_2122);
  xor g3039 (n_2130, n_3089, n_2123);
  nand g3040 (n_3090, n_2121, n_2122);
  nand g3041 (n_3091, n_2123, n_2122);
  nand g3042 (n_3092, n_2121, n_2123);
  nand g3043 (n_2158, n_3090, n_3091, n_3092);
  xor g3044 (n_3093, n_2124, n_2125);
  xor g3045 (n_2132, n_3093, n_2126);
  nand g3046 (n_3094, n_2124, n_2125);
  nand g3047 (n_3095, n_2126, n_2125);
  nand g3048 (n_3096, n_2124, n_2126);
  nand g3049 (n_2161, n_3094, n_3095, n_3096);
  xor g3050 (n_3097, n_2127, n_2128);
  xor g3051 (n_2134, n_3097, n_2129);
  nand g3052 (n_3098, n_2127, n_2128);
  nand g3053 (n_3099, n_2129, n_2128);
  nand g3054 (n_3100, n_2127, n_2129);
  nand g3055 (n_2164, n_3098, n_3099, n_3100);
  xor g3056 (n_3101, n_2130, n_2131);
  xor g3057 (n_2135, n_3101, n_2132);
  nand g3058 (n_3102, n_2130, n_2131);
  nand g3059 (n_3103, n_2132, n_2131);
  nand g3060 (n_3104, n_2130, n_2132);
  nand g3061 (n_2166, n_3102, n_3103, n_3104);
  xor g3062 (n_3105, n_2133, n_2134);
  xor g3063 (n_2137, n_3105, n_2135);
  nand g3064 (n_3106, n_2133, n_2134);
  nand g3065 (n_3107, n_2135, n_2134);
  nand g3066 (n_3108, n_2133, n_2135);
  nand g3067 (n_2168, n_3106, n_3107, n_3108);
  xor g3068 (n_3109, n_2136, n_2137);
  xor g3069 (n_176, n_3109, n_2138);
  nand g3070 (n_3110, n_2136, n_2137);
  nand g3071 (n_3111, n_2138, n_2137);
  nand g3072 (n_3112, n_2136, n_2138);
  nand g3073 (n_123, n_3110, n_3111, n_3112);
  xor g3075 (n_2156, n_3113, n_2141);
  nand g3077 (n_3115, n_2141, n_2140);
  nand g3079 (n_2181, n_3114, n_3115, n_3116);
  xor g3081 (n_2154, n_3117, n_2144);
  nand g3083 (n_3119, n_2144, n_2143);
  nand g3085 (n_2183, n_3118, n_3119, n_3120);
  xor g3086 (n_3121, n_2145, n_2146);
  xor g3087 (n_2155, n_3121, n_2147);
  nand g3088 (n_3122, n_2145, n_2146);
  nand g3089 (n_3123, n_2147, n_2146);
  nand g3090 (n_3124, n_2145, n_2147);
  nand g3091 (n_2182, n_3122, n_3123, n_3124);
  xor g3092 (n_3125, n_2148, n_2149);
  nand g3094 (n_3126, n_2148, n_2149);
  nand g3097 (n_2187, n_3126, n_3127, n_3128);
  xor g3098 (n_3129, n_2151, n_2152);
  xor g3099 (n_2160, n_3129, n_2153);
  nand g3100 (n_3130, n_2151, n_2152);
  nand g3101 (n_3131, n_2153, n_2152);
  nand g3102 (n_3132, n_2151, n_2153);
  nand g3103 (n_2188, n_3130, n_3131, n_3132);
  xor g3104 (n_3133, n_2154, n_2155);
  xor g3105 (n_2162, n_3133, n_2156);
  nand g3106 (n_3134, n_2154, n_2155);
  nand g3107 (n_3135, n_2156, n_2155);
  nand g3108 (n_3136, n_2154, n_2156);
  nand g3109 (n_2190, n_3134, n_3135, n_3136);
  xor g3110 (n_3137, n_2157, n_2158);
  xor g3111 (n_2163, n_3137, n_2159);
  nand g3112 (n_3138, n_2157, n_2158);
  nand g3113 (n_3139, n_2159, n_2158);
  nand g3114 (n_3140, n_2157, n_2159);
  nand g3115 (n_2193, n_3138, n_3139, n_3140);
  xor g3116 (n_3141, n_2160, n_2161);
  xor g3117 (n_2165, n_3141, n_2162);
  nand g3118 (n_3142, n_2160, n_2161);
  nand g3119 (n_3143, n_2162, n_2161);
  nand g3120 (n_3144, n_2160, n_2162);
  nand g3121 (n_2194, n_3142, n_3143, n_3144);
  xor g3122 (n_3145, n_2163, n_2164);
  xor g3123 (n_2167, n_3145, n_2165);
  nand g3124 (n_3146, n_2163, n_2164);
  nand g3125 (n_3147, n_2165, n_2164);
  nand g3126 (n_3148, n_2163, n_2165);
  nand g3127 (n_2197, n_3146, n_3147, n_3148);
  xor g3128 (n_3149, n_2166, n_2167);
  xor g3129 (n_175, n_3149, n_2168);
  nand g3130 (n_3150, n_2166, n_2167);
  nand g3131 (n_3151, n_2168, n_2167);
  nand g3132 (n_3152, n_2166, n_2168);
  nand g3133 (n_122, n_3150, n_3151, n_3152);
  xor g3136 (n_3153, n_2171, n_2172);
  xor g3137 (n_2185, n_3153, n_2173);
  nand g3138 (n_3154, n_2171, n_2172);
  nand g3139 (n_3155, n_2173, n_2172);
  nand g3140 (n_3156, n_2171, n_2173);
  nand g3141 (n_2209, n_3154, n_3155, n_3156);
  xor g3142 (n_3157, n_2174, n_2175);
  xor g3143 (n_2186, n_3157, n_2176);
  nand g3144 (n_3158, n_2174, n_2175);
  nand g3145 (n_3159, n_2176, n_2175);
  nand g3146 (n_3160, n_2174, n_2176);
  nand g3147 (n_2211, n_3158, n_3159, n_3160);
  xor g3148 (n_3161, n_2177, n_2178);
  xor g3149 (n_2184, n_3161, n_2179);
  nand g3150 (n_3162, n_2177, n_2178);
  nand g3151 (n_3163, n_2179, n_2178);
  nand g3152 (n_3164, n_2177, n_2179);
  nand g3153 (n_2210, n_3162, n_3163, n_3164);
  xor g3154 (n_3165, n_1521, n_2181);
  xor g3155 (n_2189, n_3165, n_2182);
  nand g3156 (n_3166, n_1521, n_2181);
  nand g3157 (n_3167, n_2182, n_2181);
  nand g3158 (n_3168, n_1521, n_2182);
  nand g3159 (n_2216, n_3166, n_3167, n_3168);
  xor g3160 (n_3169, n_2183, n_2184);
  xor g3161 (n_2191, n_3169, n_2185);
  nand g3162 (n_3170, n_2183, n_2184);
  nand g3163 (n_3171, n_2185, n_2184);
  nand g3164 (n_3172, n_2183, n_2185);
  nand g3165 (n_2217, n_3170, n_3171, n_3172);
  xor g3166 (n_3173, n_2186, n_2187);
  xor g3167 (n_2192, n_3173, n_2188);
  nand g3168 (n_3174, n_2186, n_2187);
  nand g3169 (n_3175, n_2188, n_2187);
  nand g3170 (n_3176, n_2186, n_2188);
  nand g3171 (n_2220, n_3174, n_3175, n_3176);
  xor g3172 (n_3177, n_2189, n_2190);
  xor g3173 (n_2195, n_3177, n_2191);
  nand g3174 (n_3178, n_2189, n_2190);
  nand g3175 (n_3179, n_2191, n_2190);
  nand g3176 (n_3180, n_2189, n_2191);
  nand g3177 (n_2221, n_3178, n_3179, n_3180);
  xor g3178 (n_3181, n_2192, n_2193);
  xor g3179 (n_2196, n_3181, n_2194);
  nand g3180 (n_3182, n_2192, n_2193);
  nand g3181 (n_3183, n_2194, n_2193);
  nand g3182 (n_3184, n_2192, n_2194);
  nand g3183 (n_2224, n_3182, n_3183, n_3184);
  xor g3184 (n_3185, n_2195, n_2196);
  xor g3185 (n_174, n_3185, n_2197);
  nand g3186 (n_3186, n_2195, n_2196);
  nand g3187 (n_3187, n_2197, n_2196);
  nand g3188 (n_3188, n_2195, n_2197);
  nand g3189 (n_121, n_3186, n_3187, n_3188);
  xor g3191 (n_2213, n_3189, n_2200);
  nand g3193 (n_3191, n_2200, n_2199);
  nand g3195 (n_2236, n_3190, n_3191, n_3192);
  xor g3196 (n_3193, n_2201, n_2202);
  xor g3197 (n_2214, n_3193, n_2203);
  nand g3198 (n_3194, n_2201, n_2202);
  nand g3199 (n_3195, n_2203, n_2202);
  nand g3200 (n_3196, n_2201, n_2203);
  nand g3201 (n_2238, n_3194, n_3195, n_3196);
  xor g3202 (n_3197, n_2204, n_2205);
  xor g3203 (n_2212, n_3197, n_2206);
  nand g3204 (n_3198, n_2204, n_2205);
  nand g3205 (n_3199, n_2206, n_2205);
  nand g3206 (n_3200, n_2204, n_2206);
  nand g3207 (n_2237, n_3198, n_3199, n_3200);
  xor g3209 (n_2215, n_3201, n_2209);
  nand g3213 (n_2242, n_3202, n_3203, n_3204);
  xor g3214 (n_3205, n_2210, n_2211);
  xor g3215 (n_2218, n_3205, n_2212);
  nand g3216 (n_3206, n_2210, n_2211);
  nand g3217 (n_3207, n_2212, n_2211);
  nand g3218 (n_3208, n_2210, n_2212);
  nand g3219 (n_2243, n_3206, n_3207, n_3208);
  xor g3220 (n_3209, n_2213, n_2214);
  xor g3221 (n_2219, n_3209, n_2215);
  nand g3222 (n_3210, n_2213, n_2214);
  nand g3223 (n_3211, n_2215, n_2214);
  nand g3224 (n_3212, n_2213, n_2215);
  nand g3225 (n_2246, n_3210, n_3211, n_3212);
  xor g3226 (n_3213, n_2216, n_2217);
  xor g3227 (n_2222, n_3213, n_2218);
  nand g3228 (n_3214, n_2216, n_2217);
  nand g3229 (n_3215, n_2218, n_2217);
  nand g3230 (n_3216, n_2216, n_2218);
  nand g3231 (n_2247, n_3214, n_3215, n_3216);
  xor g3232 (n_3217, n_2219, n_2220);
  xor g3233 (n_2223, n_3217, n_2221);
  nand g3234 (n_3218, n_2219, n_2220);
  nand g3235 (n_3219, n_2221, n_2220);
  nand g3236 (n_3220, n_2219, n_2221);
  nand g3237 (n_2250, n_3218, n_3219, n_3220);
  xor g3238 (n_3221, n_2222, n_2223);
  xor g3239 (n_173, n_3221, n_2224);
  nand g3240 (n_3222, n_2222, n_2223);
  nand g3241 (n_3223, n_2224, n_2223);
  nand g3242 (n_3224, n_2222, n_2224);
  nand g3243 (n_120, n_3222, n_3223, n_3224);
  xor g3246 (n_3225, n_2227, n_2228);
  xor g3247 (n_2239, n_3225, n_2229);
  nand g3248 (n_3226, n_2227, n_2228);
  nand g3249 (n_3227, n_2229, n_2228);
  nand g3250 (n_3228, n_2227, n_2229);
  nand g3251 (n_2261, n_3226, n_3227, n_3228);
  xor g3252 (n_3229, n_2230, n_2231);
  xor g3253 (n_2241, n_3229, n_2232);
  nand g3254 (n_3230, n_2230, n_2231);
  nand g3255 (n_3231, n_2232, n_2231);
  nand g3256 (n_3232, n_2230, n_2232);
  nand g3257 (n_2262, n_3230, n_3231, n_3232);
  xor g3258 (n_3233, n_2233, n_2234);
  xor g3259 (n_2240, n_3233, n_1529);
  nand g3260 (n_3234, n_2233, n_2234);
  nand g3261 (n_3235, n_1529, n_2234);
  nand g3262 (n_3236, n_2233, n_1529);
  nand g3263 (n_2265, n_3234, n_3235, n_3236);
  xor g3264 (n_3237, n_2236, n_2237);
  xor g3265 (n_2244, n_3237, n_2238);
  nand g3266 (n_3238, n_2236, n_2237);
  nand g3267 (n_3239, n_2238, n_2237);
  nand g3268 (n_3240, n_2236, n_2238);
  nand g3269 (n_2267, n_3238, n_3239, n_3240);
  xor g3270 (n_3241, n_2239, n_2240);
  xor g3271 (n_2245, n_3241, n_2241);
  nand g3272 (n_3242, n_2239, n_2240);
  nand g3273 (n_3243, n_2241, n_2240);
  nand g3274 (n_3244, n_2239, n_2241);
  nand g3275 (n_2269, n_3242, n_3243, n_3244);
  xor g3276 (n_3245, n_2242, n_2243);
  xor g3277 (n_2248, n_3245, n_2244);
  nand g3278 (n_3246, n_2242, n_2243);
  nand g3279 (n_3247, n_2244, n_2243);
  nand g3280 (n_3248, n_2242, n_2244);
  nand g3281 (n_2271, n_3246, n_3247, n_3248);
  xor g3282 (n_3249, n_2245, n_2246);
  xor g3283 (n_2249, n_3249, n_2247);
  nand g3284 (n_3250, n_2245, n_2246);
  nand g3285 (n_3251, n_2247, n_2246);
  nand g3286 (n_3252, n_2245, n_2247);
  nand g3287 (n_2274, n_3250, n_3251, n_3252);
  xor g3288 (n_3253, n_2248, n_2249);
  xor g3289 (n_172, n_3253, n_2250);
  nand g3290 (n_3254, n_2248, n_2249);
  nand g3291 (n_3255, n_2250, n_2249);
  nand g3292 (n_3256, n_2248, n_2250);
  nand g3293 (n_119, n_3254, n_3255, n_3256);
  xor g3295 (n_2264, n_3257, n_2253);
  nand g3297 (n_3259, n_2253, n_2252);
  nand g3299 (n_2286, n_3258, n_3259, n_3260);
  xor g3300 (n_3261, n_2254, n_2255);
  nand g3302 (n_3262, n_2254, n_2255);
  nand g3305 (n_2287, n_3262, n_3263, n_3264);
  xor g3306 (n_3265, n_2257, n_2258);
  xor g3307 (n_2263, n_3265, n_2259);
  nand g3308 (n_3266, n_2257, n_2258);
  nand g3309 (n_3267, n_2259, n_2258);
  nand g3310 (n_3268, n_2257, n_2259);
  nand g3311 (n_2285, n_3266, n_3267, n_3268);
  xor g3313 (n_2268, n_3269, n_2262);
  nand g3315 (n_3271, n_2262, n_2261);
  nand g3317 (n_2290, n_3270, n_3271, n_3272);
  xor g3318 (n_3273, n_2263, n_2264);
  xor g3319 (n_2270, n_3273, n_2265);
  nand g3320 (n_3274, n_2263, n_2264);
  nand g3321 (n_3275, n_2265, n_2264);
  nand g3322 (n_3276, n_2263, n_2265);
  nand g3323 (n_2293, n_3274, n_3275, n_3276);
  xor g3324 (n_3277, n_2266, n_2267);
  xor g3325 (n_2272, n_3277, n_2268);
  nand g3326 (n_3278, n_2266, n_2267);
  nand g3327 (n_3279, n_2268, n_2267);
  nand g3328 (n_3280, n_2266, n_2268);
  nand g3329 (n_2294, n_3278, n_3279, n_3280);
  xor g3330 (n_3281, n_2269, n_2270);
  xor g3331 (n_2273, n_3281, n_2271);
  nand g3332 (n_3282, n_2269, n_2270);
  nand g3333 (n_3283, n_2271, n_2270);
  nand g3334 (n_3284, n_2269, n_2271);
  nand g3335 (n_2297, n_3282, n_3283, n_3284);
  xor g3336 (n_3285, n_2272, n_2273);
  xor g3337 (n_171, n_3285, n_2274);
  nand g3338 (n_3286, n_2272, n_2273);
  nand g3339 (n_3287, n_2274, n_2273);
  nand g3340 (n_3288, n_2272, n_2274);
  nand g3341 (n_118, n_3286, n_3287, n_3288);
  xor g3344 (n_3289, n_2277, n_2278);
  xor g3345 (n_2288, n_3289, n_2279);
  nand g3346 (n_3290, n_2277, n_2278);
  nand g3347 (n_3291, n_2279, n_2278);
  nand g3348 (n_3292, n_2277, n_2279);
  nand g3349 (n_2308, n_3290, n_3291, n_3292);
  xor g3350 (n_3293, n_2280, n_2281);
  xor g3351 (n_2289, n_3293, n_2282);
  nand g3352 (n_3294, n_2280, n_2281);
  nand g3353 (n_3295, n_2282, n_2281);
  nand g3354 (n_3296, n_2280, n_2282);
  nand g3355 (n_2307, n_3294, n_3295, n_3296);
  xor g3356 (n_3297, n_2283, n_1537);
  xor g3357 (n_2291, n_3297, n_2285);
  nand g3358 (n_3298, n_2283, n_1537);
  nand g3359 (n_3299, n_2285, n_1537);
  nand g3360 (n_3300, n_2283, n_2285);
  nand g3361 (n_2312, n_3298, n_3299, n_3300);
  xor g3362 (n_3301, n_2286, n_2287);
  xor g3363 (n_2292, n_3301, n_2288);
  nand g3364 (n_3302, n_2286, n_2287);
  nand g3365 (n_3303, n_2288, n_2287);
  nand g3366 (n_3304, n_2286, n_2288);
  nand g3367 (n_2314, n_3302, n_3303, n_3304);
  xor g3368 (n_3305, n_2289, n_2290);
  xor g3369 (n_2295, n_3305, n_2291);
  nand g3370 (n_3306, n_2289, n_2290);
  nand g3371 (n_3307, n_2291, n_2290);
  nand g3372 (n_3308, n_2289, n_2291);
  nand g3373 (n_2315, n_3306, n_3307, n_3308);
  xor g3374 (n_3309, n_2292, n_2293);
  xor g3375 (n_2296, n_3309, n_2294);
  nand g3376 (n_3310, n_2292, n_2293);
  nand g3377 (n_3311, n_2294, n_2293);
  nand g3378 (n_3312, n_2292, n_2294);
  nand g3379 (n_2318, n_3310, n_3311, n_3312);
  xor g3380 (n_3313, n_2295, n_2296);
  xor g3381 (n_170, n_3313, n_2297);
  nand g3382 (n_3314, n_2295, n_2296);
  nand g3383 (n_3315, n_2297, n_2296);
  nand g3384 (n_3316, n_2295, n_2297);
  nand g3385 (n_117, n_3314, n_3315, n_3316);
  nand g3391 (n_2328, n_3318, n_3319, n_3320);
  xor g3392 (n_3321, n_2301, n_2302);
  xor g3393 (n_2311, n_3321, n_2303);
  nand g3394 (n_3322, n_2301, n_2302);
  nand g3395 (n_3323, n_2303, n_2302);
  nand g3396 (n_3324, n_2301, n_2303);
  nand g3397 (n_2329, n_3322, n_3323, n_3324);
  xor g3398 (n_3325, n_2304, n_2305);
  nand g3400 (n_3326, n_2304, n_2305);
  nand g3403 (n_2331, n_3326, n_3327, n_3328);
  xor g3404 (n_3329, n_2307, n_2308);
  xor g3405 (n_2313, n_3329, n_2309);
  nand g3406 (n_3330, n_2307, n_2308);
  nand g3407 (n_3331, n_2309, n_2308);
  nand g3408 (n_3332, n_2307, n_2309);
  nand g3409 (n_2334, n_3330, n_3331, n_3332);
  xor g3410 (n_3333, n_2310, n_2311);
  xor g3411 (n_2316, n_3333, n_2312);
  nand g3412 (n_3334, n_2310, n_2311);
  nand g3413 (n_3335, n_2312, n_2311);
  nand g3414 (n_3336, n_2310, n_2312);
  nand g3415 (n_2336, n_3334, n_3335, n_3336);
  xor g3416 (n_3337, n_2313, n_2314);
  xor g3417 (n_2317, n_3337, n_2315);
  nand g3418 (n_3338, n_2313, n_2314);
  nand g3419 (n_3339, n_2315, n_2314);
  nand g3420 (n_3340, n_2313, n_2315);
  nand g3421 (n_2338, n_3338, n_3339, n_3340);
  xor g3422 (n_3341, n_2316, n_2317);
  xor g3423 (n_169, n_3341, n_2318);
  nand g3424 (n_3342, n_2316, n_2317);
  nand g3425 (n_3343, n_2318, n_2317);
  nand g3426 (n_3344, n_2316, n_2318);
  nand g3427 (n_168, n_3342, n_3343, n_3344);
  xor g3430 (n_3345, n_2321, n_2322);
  xor g3431 (n_2332, n_3345, n_2323);
  nand g3432 (n_3346, n_2321, n_2322);
  nand g3433 (n_3347, n_2323, n_2322);
  nand g3434 (n_3348, n_2321, n_2323);
  nand g3435 (n_2347, n_3346, n_3347, n_3348);
  xor g3436 (n_3349, n_2324, n_2325);
  xor g3437 (n_2330, n_3349, n_2326);
  nand g3438 (n_3350, n_2324, n_2325);
  nand g3439 (n_3351, n_2326, n_2325);
  nand g3440 (n_3352, n_2324, n_2326);
  nand g3441 (n_2348, n_3350, n_3351, n_3352);
  xor g3442 (n_3353, n_1545, n_2328);
  xor g3443 (n_2333, n_3353, n_2329);
  nand g3444 (n_3354, n_1545, n_2328);
  nand g3445 (n_3355, n_2329, n_2328);
  nand g3446 (n_3356, n_1545, n_2329);
  nand g3447 (n_2352, n_3354, n_3355, n_3356);
  xor g3448 (n_3357, n_2330, n_2331);
  xor g3449 (n_2335, n_3357, n_2332);
  nand g3450 (n_3358, n_2330, n_2331);
  nand g3451 (n_3359, n_2332, n_2331);
  nand g3452 (n_3360, n_2330, n_2332);
  nand g3453 (n_2353, n_3358, n_3359, n_3360);
  xor g3454 (n_3361, n_2333, n_2334);
  xor g3455 (n_2337, n_3361, n_2335);
  nand g3456 (n_3362, n_2333, n_2334);
  nand g3457 (n_3363, n_2335, n_2334);
  nand g3458 (n_3364, n_2333, n_2335);
  nand g3459 (n_2356, n_3362, n_3363, n_3364);
  xor g3460 (n_3365, n_2336, n_2337);
  xor g3461 (n_116, n_3365, n_2338);
  nand g3462 (n_3366, n_2336, n_2337);
  nand g3463 (n_3367, n_2338, n_2337);
  nand g3464 (n_3368, n_2336, n_2338);
  nand g3465 (n_167, n_3366, n_3367, n_3368);
  xor g3467 (n_2350, n_3369, n_2341);
  nand g3469 (n_3371, n_2341, n_2340);
  nand g3471 (n_2366, n_3370, n_3371, n_3372);
  xor g3472 (n_3373, n_2342, n_2343);
  nand g3474 (n_3374, n_2342, n_2343);
  nand g3477 (n_2365, n_3374, n_3375, n_3376);
  xor g3479 (n_2351, n_3377, n_2347);
  nand g3482 (n_3380, n_2345, n_2347);
  nand g3483 (n_2369, n_3378, n_3379, n_3380);
  xor g3484 (n_3381, n_2348, n_2349);
  xor g3485 (n_2354, n_3381, n_2350);
  nand g3486 (n_3382, n_2348, n_2349);
  nand g3487 (n_3383, n_2350, n_2349);
  nand g3488 (n_3384, n_2348, n_2350);
  nand g3489 (n_2370, n_3382, n_3383, n_3384);
  xor g3490 (n_3385, n_2351, n_2352);
  xor g3491 (n_2355, n_3385, n_2353);
  nand g3492 (n_3386, n_2351, n_2352);
  nand g3493 (n_3387, n_2353, n_2352);
  nand g3494 (n_3388, n_2351, n_2353);
  nand g3495 (n_2373, n_3386, n_3387, n_3388);
  xor g3496 (n_3389, n_2354, n_2355);
  xor g3497 (n_115, n_3389, n_2356);
  nand g3498 (n_3390, n_2354, n_2355);
  nand g3499 (n_3391, n_2356, n_2355);
  nand g3500 (n_3392, n_2354, n_2356);
  nand g3501 (n_114, n_3390, n_3391, n_3392);
  xor g3504 (n_3393, n_2359, n_2360);
  xor g3505 (n_2367, n_3393, n_2361);
  nand g3506 (n_3394, n_2359, n_2360);
  nand g3507 (n_3395, n_2361, n_2360);
  nand g3508 (n_3396, n_2359, n_2361);
  nand g3509 (n_2381, n_3394, n_3395, n_3396);
  xor g3510 (n_3397, n_2362, n_2363);
  xor g3511 (n_2368, n_3397, n_1553);
  nand g3512 (n_3398, n_2362, n_2363);
  nand g3513 (n_3399, n_1553, n_2363);
  nand g3514 (n_3400, n_2362, n_1553);
  nand g3515 (n_2383, n_3398, n_3399, n_3400);
  xor g3516 (n_3401, n_2365, n_2366);
  xor g3517 (n_2371, n_3401, n_2367);
  nand g3518 (n_3402, n_2365, n_2366);
  nand g3519 (n_3403, n_2367, n_2366);
  nand g3520 (n_3404, n_2365, n_2367);
  nand g3521 (n_2386, n_3402, n_3403, n_3404);
  xor g3522 (n_3405, n_2368, n_2369);
  xor g3523 (n_2372, n_3405, n_2370);
  nand g3524 (n_3406, n_2368, n_2369);
  nand g3525 (n_3407, n_2370, n_2369);
  nand g3526 (n_3408, n_2368, n_2370);
  nand g3527 (n_2388, n_3406, n_3407, n_3408);
  xor g3528 (n_3409, n_2371, n_2372);
  xor g3529 (n_166, n_3409, n_2373);
  nand g3530 (n_3410, n_2371, n_2372);
  nand g3531 (n_3411, n_2373, n_2372);
  nand g3532 (n_3412, n_2371, n_2373);
  nand g3533 (n_113, n_3410, n_3411, n_3412);
  nand g3539 (n_2396, n_3414, n_3415, n_3416);
  xor g3540 (n_3417, n_2377, n_2378);
  xor g3541 (n_2382, n_3417, n_2379);
  nand g3542 (n_3418, n_2377, n_2378);
  nand g3543 (n_3419, n_2379, n_2378);
  nand g3544 (n_3420, n_2377, n_2379);
  nand g3545 (n_2397, n_3418, n_3419, n_3420);
  xor g3547 (n_2385, n_3421, n_2382);
  nand g3549 (n_3423, n_2382, n_2381);
  nand g3551 (n_2400, n_3422, n_3423, n_3424);
  xor g3552 (n_3425, n_2383, n_2384);
  xor g3553 (n_2387, n_3425, n_2385);
  nand g3554 (n_3426, n_2383, n_2384);
  nand g3555 (n_3427, n_2385, n_2384);
  nand g3556 (n_3428, n_2383, n_2385);
  nand g3557 (n_2402, n_3426, n_3427, n_3428);
  xor g3558 (n_3429, n_2386, n_2387);
  xor g3559 (n_165, n_3429, n_2388);
  nand g3560 (n_3430, n_2386, n_2387);
  nand g3561 (n_3431, n_2388, n_2387);
  nand g3562 (n_3432, n_2386, n_2388);
  nand g3563 (n_112, n_3430, n_3431, n_3432);
  xor g3566 (n_3433, n_2391, n_2392);
  xor g3567 (n_2398, n_3433, n_2393);
  nand g3568 (n_3434, n_2391, n_2392);
  nand g3569 (n_3435, n_2393, n_2392);
  nand g3570 (n_3436, n_2391, n_2393);
  nand g3571 (n_2409, n_3434, n_3435, n_3436);
  xor g3572 (n_3437, n_2394, n_1561);
  xor g3573 (n_2399, n_3437, n_2396);
  nand g3574 (n_3438, n_2394, n_1561);
  nand g3575 (n_3439, n_2396, n_1561);
  nand g3576 (n_3440, n_2394, n_2396);
  nand g3577 (n_2412, n_3438, n_3439, n_3440);
  xor g3578 (n_3441, n_2397, n_2398);
  xor g3579 (n_2401, n_3441, n_2399);
  nand g3580 (n_3442, n_2397, n_2398);
  nand g3581 (n_3443, n_2399, n_2398);
  nand g3582 (n_3444, n_2397, n_2399);
  nand g3583 (n_2414, n_3442, n_3443, n_3444);
  xor g3584 (n_3445, n_2400, n_2401);
  xor g3585 (n_164, n_3445, n_2402);
  nand g3586 (n_3446, n_2400, n_2401);
  nand g3587 (n_3447, n_2402, n_2401);
  nand g3588 (n_3448, n_2400, n_2402);
  nand g3589 (n_163, n_3446, n_3447, n_3448);
  nand g3595 (n_2421, n_3450, n_3451, n_3452);
  xor g3596 (n_3453, n_2406, n_2407);
  nand g3598 (n_3454, n_2406, n_2407);
  nand g3601 (n_2423, n_3454, n_3455, n_3456);
  xor g3602 (n_3457, n_2409, n_2410);
  xor g3603 (n_2413, n_3457, n_2411);
  nand g3604 (n_3458, n_2409, n_2410);
  nand g3605 (n_3459, n_2411, n_2410);
  nand g3606 (n_3460, n_2409, n_2411);
  nand g3607 (n_2425, n_3458, n_3459, n_3460);
  xor g3608 (n_3461, n_2412, n_2413);
  xor g3609 (n_111, n_3461, n_2414);
  nand g3610 (n_3462, n_2412, n_2413);
  nand g3611 (n_3463, n_2414, n_2413);
  nand g3612 (n_3464, n_2412, n_2414);
  nand g3613 (n_162, n_3462, n_3463, n_3464);
  xor g3616 (n_3465, n_2417, n_2418);
  xor g3617 (n_2422, n_3465, n_2419);
  nand g3618 (n_3466, n_2417, n_2418);
  nand g3619 (n_3467, n_2419, n_2418);
  nand g3620 (n_3468, n_2417, n_2419);
  nand g3621 (n_2431, n_3466, n_3467, n_3468);
  xor g3622 (n_3469, n_1569, n_2421);
  xor g3623 (n_2424, n_3469, n_2422);
  nand g3624 (n_3470, n_1569, n_2421);
  nand g3625 (n_3471, n_2422, n_2421);
  nand g3626 (n_3472, n_1569, n_2422);
  nand g3627 (n_2434, n_3470, n_3471, n_3472);
  xor g3628 (n_3473, n_2423, n_2424);
  xor g3629 (n_110, n_3473, n_2425);
  nand g3630 (n_3474, n_2423, n_2424);
  nand g3631 (n_3475, n_2425, n_2424);
  nand g3632 (n_3476, n_2423, n_2425);
  nand g3633 (n_109, n_3474, n_3475, n_3476);
  xor g3635 (n_2432, n_3477, n_2428);
  nand g3637 (n_3479, n_2428, n_2427);
  nand g3639 (n_2440, n_3478, n_3479, n_3480);
  xor g3641 (n_2433, n_3481, n_2431);
  nand g3645 (n_2442, n_3482, n_3483, n_3484);
  xor g3646 (n_3485, n_2432, n_2433);
  xor g3647 (n_161, n_3485, n_2434);
  nand g3648 (n_3486, n_2432, n_2433);
  nand g3649 (n_3487, n_2434, n_2433);
  nand g3650 (n_3488, n_2432, n_2434);
  nand g3651 (n_160, n_3486, n_3487, n_3488);
  xor g3654 (n_3489, n_2437, n_2438);
  xor g3655 (n_2441, n_3489, n_1577);
  nand g3656 (n_3490, n_2437, n_2438);
  nand g3657 (n_3491, n_1577, n_2438);
  nand g3658 (n_3492, n_2437, n_1577);
  nand g3659 (n_2448, n_3490, n_3491, n_3492);
  xor g3660 (n_3493, n_2440, n_2441);
  xor g3661 (n_108, n_3493, n_2442);
  nand g3662 (n_3494, n_2440, n_2441);
  nand g3663 (n_3495, n_2442, n_2441);
  nand g3664 (n_3496, n_2440, n_2442);
  nand g3665 (n_159, n_3494, n_3495, n_3496);
  xor g3667 (n_2447, n_3497, n_2445);
  nand g3671 (n_2453, n_3498, n_3499, n_3500);
  xor g3673 (n_107, n_3501, n_2448);
  nand g3675 (n_3503, n_2448, n_2447);
  nand g3677 (n_158, n_3502, n_3503, n_3504);
  xor g3680 (n_3505, n_2451, n_1585);
  xor g3681 (n_106, n_3505, n_2453);
  nand g3682 (n_3506, n_2451, n_1585);
  nand g3683 (n_3507, n_2453, n_1585);
  nand g3684 (n_3508, n_2451, n_2453);
  nand g3685 (n_157, n_3506, n_3507, n_3508);
  nor g3705 (n_3535, n_152, n_204);
  nand g3706 (n_3530, n_152, n_204);
  nor g3709 (n_3541, n_150, n_202);
  nand g3710 (n_3536, n_150, n_202);
  nor g3711 (n_3537, n_149, n_201);
  nand g3712 (n_3538, n_149, n_201);
  nor g3713 (n_3547, n_148, n_200);
  nand g3714 (n_3542, n_148, n_200);
  nor g3715 (n_3543, n_147, n_199);
  nand g3716 (n_3544, n_147, n_199);
  nor g3717 (n_3553, n_146, n_198);
  nand g3718 (n_3548, n_146, n_198);
  nor g3719 (n_3549, n_145, n_197);
  nand g3720 (n_3550, n_145, n_197);
  nor g3721 (n_3559, n_144, n_196);
  nand g3722 (n_3554, n_144, n_196);
  nor g3723 (n_3555, n_143, n_195);
  nand g3724 (n_3556, n_143, n_195);
  nor g3725 (n_3565, n_142, n_194);
  nand g3726 (n_3560, n_142, n_194);
  nor g3727 (n_3561, n_141, n_193);
  nand g3728 (n_3562, n_141, n_193);
  nor g3729 (n_3571, n_140, n_192);
  nand g3730 (n_3566, n_140, n_192);
  nor g3731 (n_3567, n_139, n_191);
  nand g3732 (n_3568, n_139, n_191);
  nor g3733 (n_3577, n_138, n_190);
  nand g3734 (n_3572, n_138, n_190);
  nor g3735 (n_3573, n_137, n_189);
  nand g3736 (n_3574, n_137, n_189);
  nor g3737 (n_3583, n_136, n_188);
  nand g3738 (n_3578, n_136, n_188);
  nor g3739 (n_3579, n_135, n_187);
  nand g3740 (n_3580, n_135, n_187);
  nor g3741 (n_3589, n_134, n_186);
  nand g3742 (n_3584, n_134, n_186);
  nor g3743 (n_3585, n_133, n_185);
  nand g3744 (n_3586, n_133, n_185);
  nor g3745 (n_3595, n_132, n_184);
  nand g3746 (n_3590, n_132, n_184);
  nor g3747 (n_3591, n_131, n_183);
  nand g3748 (n_3592, n_131, n_183);
  nor g3749 (n_3601, n_130, n_182);
  nand g3750 (n_3596, n_130, n_182);
  nor g3751 (n_3597, n_129, n_181);
  nand g3752 (n_3598, n_129, n_181);
  nor g3753 (n_3607, n_128, n_180);
  nand g3754 (n_3602, n_128, n_180);
  nor g3755 (n_3603, n_127, n_179);
  nand g3756 (n_3604, n_127, n_179);
  nor g3757 (n_3613, n_126, n_178);
  nand g3758 (n_3608, n_126, n_178);
  nor g3759 (n_3609, n_125, n_177);
  nand g3760 (n_3610, n_125, n_177);
  nor g3761 (n_3619, n_124, n_176);
  nand g3762 (n_3614, n_124, n_176);
  nor g3763 (n_3615, n_123, n_175);
  nand g3764 (n_3616, n_123, n_175);
  nor g3765 (n_3625, n_122, n_174);
  nand g3766 (n_3620, n_122, n_174);
  nor g3767 (n_3621, n_121, n_173);
  nand g3768 (n_3622, n_121, n_173);
  nor g3769 (n_3631, n_120, n_172);
  nand g3770 (n_3626, n_120, n_172);
  nor g3771 (n_3627, n_119, n_171);
  nand g3772 (n_3628, n_119, n_171);
  nor g3773 (n_3637, n_118, n_170);
  nand g3774 (n_3632, n_118, n_170);
  nor g3775 (n_3633, n_117, n_169);
  nand g3776 (n_3634, n_117, n_169);
  nor g3777 (n_3643, n_116, n_168);
  nand g3778 (n_3638, n_116, n_168);
  nor g3779 (n_3639, n_115, n_167);
  nand g3780 (n_3640, n_115, n_167);
  nor g3781 (n_3649, n_114, n_166);
  nand g3782 (n_3644, n_114, n_166);
  nor g3783 (n_3645, n_113, n_165);
  nand g3784 (n_3646, n_113, n_165);
  nor g3785 (n_3655, n_112, n_164);
  nand g3786 (n_3650, n_112, n_164);
  nor g3787 (n_3651, n_111, n_163);
  nand g3788 (n_3652, n_111, n_163);
  nor g3789 (n_3661, n_110, n_162);
  nand g3790 (n_3656, n_110, n_162);
  nor g3791 (n_3657, n_109, n_161);
  nand g3792 (n_3658, n_109, n_161);
  nor g3793 (n_3667, n_108, n_160);
  nand g3794 (n_3662, n_108, n_160);
  nor g3795 (n_3663, n_107, n_159);
  nand g3796 (n_3664, n_107, n_159);
  nor g3797 (n_3671, n_106, n_158);
  nand g3798 (n_3668, n_106, n_158);
  nor g3812 (n_3539, n_3536, n_3537);
  nor g3815 (n_3683, n_3541, n_3537);
  nor g3816 (n_3545, n_3542, n_3543);
  nor g3819 (n_3691, n_3547, n_3543);
  nor g3820 (n_3551, n_3548, n_3549);
  nor g3823 (n_3693, n_3553, n_3549);
  nor g3824 (n_3557, n_3554, n_3555);
  nor g3827 (n_3701, n_3559, n_3555);
  nor g3828 (n_3563, n_3560, n_3561);
  nor g3831 (n_3703, n_3565, n_3561);
  nor g3832 (n_3569, n_3566, n_3567);
  nor g3835 (n_3711, n_3571, n_3567);
  nor g3836 (n_3575, n_3572, n_3573);
  nor g3839 (n_3713, n_3577, n_3573);
  nor g3840 (n_3581, n_3578, n_3579);
  nor g3843 (n_3721, n_3583, n_3579);
  nor g3844 (n_3587, n_3584, n_3585);
  nor g3847 (n_3723, n_3589, n_3585);
  nor g3848 (n_3593, n_3590, n_3591);
  nor g3851 (n_3731, n_3595, n_3591);
  nor g3852 (n_3599, n_3596, n_3597);
  nor g3855 (n_3733, n_3601, n_3597);
  nor g3856 (n_3605, n_3602, n_3603);
  nor g3859 (n_3741, n_3607, n_3603);
  nor g3860 (n_3611, n_3608, n_3609);
  nor g3863 (n_3743, n_3613, n_3609);
  nor g3864 (n_3617, n_3614, n_3615);
  nor g3867 (n_3751, n_3619, n_3615);
  nor g3868 (n_3623, n_3620, n_3621);
  nor g3871 (n_3753, n_3625, n_3621);
  nor g3872 (n_3629, n_3626, n_3627);
  nor g3875 (n_3761, n_3631, n_3627);
  nor g3876 (n_3635, n_3632, n_3633);
  nor g3879 (n_3763, n_3637, n_3633);
  nor g3880 (n_3641, n_3638, n_3639);
  nor g3883 (n_3771, n_3643, n_3639);
  nor g3884 (n_3647, n_3644, n_3645);
  nor g3887 (n_3773, n_3649, n_3645);
  nor g3888 (n_3653, n_3650, n_3651);
  nor g3891 (n_3781, n_3655, n_3651);
  nor g3892 (n_3659, n_3656, n_3657);
  nor g3895 (n_3783, n_3661, n_3657);
  nor g3896 (n_3665, n_3662, n_3663);
  nor g3899 (n_3791, n_3667, n_3663);
  nor g3915 (n_3689, n_3553, n_3688);
  nand g3924 (n_3808, n_3691, n_3693);
  nor g3925 (n_3699, n_3565, n_3698);
  nand g3934 (n_3816, n_3701, n_3703);
  nor g3935 (n_3709, n_3577, n_3708);
  nand g3944 (n_3823, n_3711, n_3713);
  nor g3945 (n_3719, n_3589, n_3718);
  nand g3954 (n_3831, n_3721, n_3723);
  nor g3955 (n_3729, n_3601, n_3728);
  nand g3964 (n_3838, n_3731, n_3733);
  nor g3965 (n_3739, n_3613, n_3738);
  nand g3974 (n_3846, n_3741, n_3743);
  nor g3975 (n_3749, n_3625, n_3748);
  nand g3984 (n_3853, n_3751, n_3753);
  nor g3985 (n_3759, n_3637, n_3758);
  nand g3994 (n_3861, n_3761, n_3763);
  nor g3995 (n_3769, n_3649, n_3768);
  nand g4004 (n_3868, n_3771, n_3773);
  nor g4005 (n_3779, n_3661, n_3778);
  nand g4014 (n_3876, n_3781, n_3783);
  nor g4015 (n_3789, n_3671, n_3788);
  nor g4031 (n_3806, n_3559, n_3805);
  nor g4034 (n_3890, n_3559, n_3808);
  nor g4040 (n_3814, n_3812, n_3805);
  nor g4043 (n_3896, n_3808, n_3812);
  nor g4044 (n_3818, n_3816, n_3805);
  nor g4047 (n_3899, n_3808, n_3816);
  nor g4048 (n_3821, n_3583, n_3820);
  nor g4051 (n_3984, n_3583, n_3823);
  nor g4057 (n_3829, n_3827, n_3820);
  nor g4060 (n_3990, n_3823, n_3827);
  nor g4061 (n_3833, n_3831, n_3820);
  nor g4064 (n_3905, n_3823, n_3831);
  nor g4065 (n_3836, n_3607, n_3835);
  nor g4068 (n_3918, n_3607, n_3838);
  nor g4074 (n_3844, n_3842, n_3835);
  nor g4077 (n_3928, n_3838, n_3842);
  nor g4078 (n_3848, n_3846, n_3835);
  nor g4081 (n_3933, n_3838, n_3846);
  nor g4082 (n_3851, n_3631, n_3850);
  nor g4085 (n_4047, n_3631, n_3853);
  nor g4091 (n_3859, n_3857, n_3850);
  nor g4094 (n_4053, n_3853, n_3857);
  nor g4095 (n_3863, n_3861, n_3850);
  nor g4098 (n_3941, n_3853, n_3861);
  nor g4099 (n_3866, n_3655, n_3865);
  nor g4102 (n_3954, n_3655, n_3868);
  nor g4108 (n_3874, n_3872, n_3865);
  nor g4111 (n_3964, n_3868, n_3872);
  nor g4112 (n_3878, n_3876, n_3865);
  nor g4115 (n_3969, n_3868, n_3876);
  nand g4118 (n_4112, n_3542, n_3882);
  nand g4120 (n_4114, n_3688, n_3883);
  nand g4123 (n_4117, n_3886, n_3887);
  nand g4126 (n_4120, n_3805, n_3889);
  nand g4128 (n_4123, n_3891, n_3892);
  nand g4130 (n_4125, n_3894, n_3895);
  nand g4132 (n_4128, n_3897, n_3898);
  nand g4134 (n_3974, n_3900, n_3901);
  nor g4135 (n_3903, n_3595, n_3902);
  nand g4144 (n_3998, n_3731, n_3905);
  nor g4145 (n_3912, n_3910, n_3902);
  nor g4150 (n_3915, n_3838, n_3902);
  nand g4159 (n_4010, n_3905, n_3918);
  nand g4164 (n_4014, n_3905, n_3923);
  nand g4169 (n_4018, n_3905, n_3928);
  nand g4174 (n_4022, n_3905, n_3933);
  nor g4175 (n_3939, n_3643, n_3938);
  nand g4184 (n_4061, n_3771, n_3941);
  nor g4185 (n_3948, n_3946, n_3938);
  nor g4190 (n_3951, n_3868, n_3938);
  nand g4199 (n_4073, n_3941, n_3954);
  nand g4204 (n_4077, n_3941, n_3959);
  nand g4209 (n_4081, n_3941, n_3964);
  nand g4214 (n_4029, n_3941, n_3969);
  nand g4217 (n_4132, n_3566, n_3976);
  nand g4218 (n_3977, n_3711, n_3974);
  nand g4219 (n_4134, n_3708, n_3977);
  nand g4222 (n_4137, n_3980, n_3981);
  nand g4225 (n_4140, n_3820, n_3983);
  nand g4226 (n_3986, n_3984, n_3974);
  nand g4227 (n_4143, n_3985, n_3986);
  nand g4228 (n_3989, n_3987, n_3974);
  nand g4229 (n_4145, n_3988, n_3989);
  nand g4230 (n_3992, n_3990, n_3974);
  nand g4231 (n_4148, n_3991, n_3992);
  nand g4232 (n_3993, n_3905, n_3974);
  nand g4233 (n_4150, n_3902, n_3993);
  nand g4236 (n_4153, n_3996, n_3997);
  nand g4239 (n_4155, n_4000, n_4001);
  nand g4242 (n_4158, n_4004, n_4005);
  nand g4245 (n_4161, n_4008, n_4009);
  nand g4248 (n_4164, n_4012, n_4013);
  nand g4251 (n_4166, n_4016, n_4017);
  nand g4254 (n_4169, n_4020, n_4021);
  nand g4257 (n_4037, n_4024, n_4025);
  nor g4258 (n_4027, n_3667, n_4026);
  nor g4261 (n_4087, n_3667, n_4029);
  nor g4267 (n_4035, n_4033, n_4026);
  nor g4270 (n_4093, n_4033, n_4029);
  nand g4273 (n_4173, n_3614, n_4039);
  nand g4274 (n_4040, n_3751, n_4037);
  nand g4275 (n_4175, n_3748, n_4040);
  nand g4278 (n_4178, n_4043, n_4044);
  nand g4281 (n_4181, n_3850, n_4046);
  nand g4282 (n_4049, n_4047, n_4037);
  nand g4283 (n_4184, n_4048, n_4049);
  nand g4284 (n_4052, n_4050, n_4037);
  nand g4285 (n_4186, n_4051, n_4052);
  nand g4286 (n_4055, n_4053, n_4037);
  nand g4287 (n_4189, n_4054, n_4055);
  nand g4288 (n_4056, n_3941, n_4037);
  nand g4289 (n_4191, n_3938, n_4056);
  nand g4292 (n_4194, n_4059, n_4060);
  nand g4295 (n_4196, n_4063, n_4064);
  nand g4298 (n_4199, n_4067, n_4068);
  nand g4301 (n_4202, n_4071, n_4072);
  nand g4304 (n_4205, n_4075, n_4076);
  nand g4307 (n_4207, n_4079, n_4080);
  nand g4310 (n_4210, n_4083, n_4084);
  nand g4313 (n_4213, n_4026, n_4086);
  nand g4314 (n_4089, n_4087, n_4037);
  nand g4315 (n_4216, n_4088, n_4089);
  nand g4316 (n_4092, n_4090, n_4037);
  nand g4317 (n_4218, n_4091, n_4092);
  nand g4318 (n_4095, n_4093, n_4037);
  nand g4319 (n_4221, n_4094, n_4095);
  xnor g4333 (Z[6], n_3533, n_4106);
  xnor g4341 (Z[9], n_4112, n_4113);
  xnor g4343 (Z[10], n_4114, n_4115);
  xnor g4346 (Z[11], n_4117, n_4118);
  xnor g4349 (Z[12], n_4120, n_4121);
  xnor g4352 (Z[13], n_4123, n_4124);
  xnor g4354 (Z[14], n_4125, n_4126);
  xnor g4357 (Z[15], n_4128, n_4129);
  xnor g4359 (Z[16], n_3974, n_4130);
  xnor g4362 (Z[17], n_4132, n_4133);
  xnor g4364 (Z[18], n_4134, n_4135);
  xnor g4367 (Z[19], n_4137, n_4138);
  xnor g4370 (Z[20], n_4140, n_4141);
  xnor g4373 (Z[21], n_4143, n_4144);
  xnor g4375 (Z[22], n_4145, n_4146);
  xnor g4378 (Z[23], n_4148, n_4149);
  xnor g4380 (Z[24], n_4150, n_4151);
  xnor g4383 (Z[25], n_4153, n_4154);
  xnor g4385 (Z[26], n_4155, n_4156);
  xnor g4388 (Z[27], n_4158, n_4159);
  xnor g4391 (Z[28], n_4161, n_4162);
  xnor g4394 (Z[29], n_4164, n_4165);
  xnor g4396 (Z[30], n_4166, n_4167);
  xnor g4399 (Z[31], n_4169, n_4170);
  xnor g4401 (Z[32], n_4037, n_4171);
  xnor g4404 (Z[33], n_4173, n_4174);
  xnor g4406 (Z[34], n_4175, n_4176);
  xnor g4409 (Z[35], n_4178, n_4179);
  xnor g4412 (Z[36], n_4181, n_4182);
  xnor g4415 (Z[37], n_4184, n_4185);
  xnor g4417 (Z[38], n_4186, n_4187);
  xnor g4420 (Z[39], n_4189, n_4190);
  xnor g4422 (Z[40], n_4191, n_4192);
  xnor g4425 (Z[41], n_4194, n_4195);
  xnor g4427 (Z[42], n_4196, n_4197);
  xnor g4430 (Z[43], n_4199, n_4200);
  xnor g4433 (Z[44], n_4202, n_4203);
  xnor g4436 (Z[45], n_4205, n_4206);
  xnor g4438 (Z[46], n_4207, n_4208);
  xnor g4441 (Z[47], n_4210, n_4211);
  xnor g4444 (Z[48], n_4213, n_4214);
  xnor g4447 (Z[49], n_4216, n_4217);
  xnor g4449 (Z[50], n_4218, n_4219);
  xnor g4452 (Z[51], n_4221, n_4222);
  and g4454 (n_405, wc, n_404);
  not gc (wc, A[0]);
  and g4455 (n_502, wc0, n_501);
  not gc0 (wc0, A[0]);
  and g4456 (n_599, wc1, n_598);
  not gc1 (wc1, A[0]);
  and g4457 (n_696, wc2, n_695);
  not gc2 (wc2, A[0]);
  and g4458 (n_793, wc3, n_792);
  not gc3 (wc3, A[0]);
  and g4459 (n_890, wc4, n_889);
  not gc4 (wc4, A[0]);
  and g4460 (n_987, wc5, n_986);
  not gc5 (wc5, A[0]);
  and g4461 (n_1084, wc6, n_1083);
  not gc6 (wc6, A[0]);
  and g4462 (n_1181, wc7, n_1180);
  not gc7 (wc7, A[0]);
  and g4463 (n_1278, wc8, n_1277);
  not gc8 (wc8, A[0]);
  and g4464 (n_1375, wc9, n_1374);
  not gc9 (wc9, A[0]);
  and g4465 (n_1472, wc10, n_1471);
  not gc10 (wc10, A[0]);
  and g4466 (n_315, n_313, wc11);
  not gc11 (wc11, n_311);
  and g4467 (n_412, n_410, wc12);
  not gc12 (wc12, n_408);
  and g4468 (n_509, n_507, wc13);
  not gc13 (wc13, n_505);
  and g4469 (n_606, n_604, wc14);
  not gc14 (wc14, n_602);
  and g4470 (n_703, n_701, wc15);
  not gc15 (wc15, n_699);
  and g4471 (n_800, n_798, wc16);
  not gc16 (wc16, n_796);
  and g4472 (n_897, n_895, wc17);
  not gc17 (wc17, n_893);
  and g4473 (n_994, n_992, wc18);
  not gc18 (wc18, n_990);
  and g4474 (n_1091, n_1089, wc19);
  not gc19 (wc19, n_1087);
  and g4475 (n_1188, n_1186, wc20);
  not gc20 (wc20, n_1184);
  and g4476 (n_1285, n_1283, wc21);
  not gc21 (wc21, n_1281);
  and g4477 (n_1382, n_1380, wc22);
  not gc22 (wc22, n_1378);
  xnor g4501 (n_2897, n_1972, n_1497);
  or g4502 (n_2898, n_1497, wc23);
  not gc23 (wc23, n_1972);
  or g4503 (n_2900, n_1497, wc24);
  not gc24 (wc24, n_1973);
  xnor g4504 (n_3029, n_2075, n_1509);
  or g4505 (n_3030, n_1509, wc25);
  not gc25 (wc25, n_2075);
  or g4506 (n_3032, n_1509, wc26);
  not gc26 (wc26, n_2076);
  xnor g4507 (n_3113, n_2140, n_1517);
  or g4508 (n_3114, n_1517, wc27);
  not gc27 (wc27, n_2140);
  or g4509 (n_3116, n_1517, wc28);
  not gc28 (wc28, n_2141);
  xnor g4510 (n_3189, n_2199, n_1525);
  or g4511 (n_3190, n_1525, wc29);
  not gc29 (wc29, n_2199);
  or g4512 (n_3192, n_1525, wc30);
  not gc30 (wc30, n_2200);
  xnor g4513 (n_3257, n_2252, n_1533);
  or g4514 (n_3258, n_1533, wc31);
  not gc31 (wc31, n_2252);
  or g4515 (n_3260, n_1533, wc32);
  not gc32 (wc32, n_2253);
  xnor g4516 (n_3317, n_2299, n_1541);
  or g4517 (n_3318, n_1541, wc33);
  not gc33 (wc33, n_2299);
  xnor g4518 (n_3369, n_2340, n_1549);
  or g4519 (n_3370, n_1549, wc34);
  not gc34 (wc34, n_2340);
  or g4520 (n_3372, n_1549, wc35);
  not gc35 (wc35, n_2341);
  xnor g4521 (n_3413, n_2375, n_1557);
  or g4522 (n_3414, n_1557, wc36);
  not gc36 (wc36, n_2375);
  xnor g4523 (n_3449, n_2404, n_1565);
  or g4524 (n_3450, n_1565, wc37);
  not gc37 (wc37, n_2404);
  xnor g4525 (n_3477, n_2427, n_1573);
  or g4526 (n_3478, n_1573, wc38);
  not gc38 (wc38, n_2427);
  or g4527 (n_3480, n_1573, wc39);
  not gc39 (wc39, n_2428);
  or g4528 (n_3500, n_1581, wc40);
  not gc40 (wc40, n_2445);
  xnor g4530 (n_2949, n_402, n_2013);
  or g4531 (n_2950, wc41, n_402);
  not gc41 (wc41, n_2013);
  or g4532 (n_2952, wc42, n_402);
  not gc42 (wc42, n_2014);
  xnor g4533 (n_3033, n_499, n_2078);
  or g4534 (n_3034, wc43, n_499);
  not gc43 (wc43, n_2078);
  or g4535 (n_3036, wc44, n_499);
  not gc44 (wc44, n_2079);
  xnor g4536 (n_3117, n_596, n_2143);
  or g4537 (n_3118, wc45, n_596);
  not gc45 (wc45, n_2143);
  or g4538 (n_3120, wc46, n_596);
  not gc46 (wc46, n_2144);
  xnor g4539 (n_2157, n_1513, n_3125);
  or g4540 (n_3127, n_1513, wc47);
  not gc47 (wc47, n_2149);
  or g4541 (n_3128, n_1513, wc48);
  not gc48 (wc48, n_2148);
  xor g4542 (n_3201, n_693, n_1521);
  or g4543 (n_3202, n_693, n_1521);
  xnor g4544 (n_2266, n_790, n_3261);
  or g4545 (n_3263, wc49, n_790);
  not gc49 (wc49, n_2255);
  or g4546 (n_3264, wc50, n_790);
  not gc50 (wc50, n_2254);
  xnor g4547 (n_2309, n_887, n_3317);
  or g4548 (n_3319, wc51, n_887);
  not gc51 (wc51, n_2299);
  or g4549 (n_3320, n_887, n_1541);
  xnor g4550 (n_2310, n_1537, n_3325);
  or g4551 (n_3327, n_1537, wc52);
  not gc52 (wc52, n_2305);
  or g4552 (n_3328, n_1537, wc53);
  not gc53 (wc53, n_2304);
  xnor g4553 (n_2349, n_984, n_3373);
  or g4554 (n_3375, wc54, n_984);
  not gc54 (wc54, n_2343);
  or g4555 (n_3376, wc55, n_984);
  not gc55 (wc55, n_2342);
  xnor g4556 (n_3377, n_2345, n_1545);
  or g4557 (n_3378, n_1545, wc56);
  not gc56 (wc56, n_2345);
  xnor g4558 (n_2384, n_1081, n_3413);
  or g4559 (n_3415, wc57, n_1081);
  not gc57 (wc57, n_2375);
  or g4560 (n_3416, n_1081, n_1557);
  xnor g4561 (n_2410, n_1178, n_3449);
  or g4562 (n_3451, wc58, n_1178);
  not gc58 (wc58, n_2404);
  or g4563 (n_3452, n_1178, n_1565);
  xnor g4564 (n_2411, n_1561, n_3453);
  or g4565 (n_3455, n_1561, wc59);
  not gc59 (wc59, n_2407);
  or g4566 (n_3456, n_1561, wc60);
  not gc60 (wc60, n_2406);
  xor g4567 (n_3481, n_1275, n_1569);
  or g4568 (n_3482, n_1275, n_1569);
  xor g4569 (n_3497, n_1372, n_1581);
  or g4570 (n_3498, n_1372, n_1581);
  or g4571 (n_3499, wc61, n_1372);
  not gc61 (wc61, n_2445);
  and g4572 (n_3533, wc62, n_151);
  not gc62 (wc62, n_3530);
  xnor g4574 (n_3001, n_1501, n_2054);
  or g4575 (n_3002, wc63, n_1501);
  not gc63 (wc63, n_2054);
  or g4576 (n_3004, wc64, n_1501);
  not gc64 (wc64, n_2055);
  xnor g4577 (n_3045, n_1505, n_2087);
  or g4578 (n_3046, wc65, n_1505);
  not gc65 (wc65, n_2087);
  or g4579 (n_3048, wc66, n_1505);
  not gc66 (wc66, n_2088);
  or g4580 (n_3203, wc67, n_1521);
  not gc67 (wc67, n_2209);
  or g4581 (n_3204, wc68, n_693);
  not gc68 (wc68, n_2209);
  xnor g4582 (n_3269, n_1529, n_2261);
  or g4583 (n_3270, wc69, n_1529);
  not gc69 (wc69, n_2261);
  or g4584 (n_3272, wc70, n_1529);
  not gc70 (wc70, n_2262);
  or g4585 (n_3379, wc71, n_1545);
  not gc71 (wc71, n_2347);
  xnor g4586 (n_3421, n_1553, n_2381);
  or g4587 (n_3422, wc72, n_1553);
  not gc72 (wc72, n_2381);
  or g4588 (n_3424, wc73, n_1553);
  not gc73 (wc73, n_2382);
  or g4589 (n_3483, wc74, n_1569);
  not gc74 (wc74, n_2431);
  or g4590 (n_3484, wc75, n_1275);
  not gc75 (wc75, n_2431);
  xnor g4591 (n_105, n_1469, n_1585);
  or g4593 (n_4101, wc76, n_3535);
  not gc76 (wc76, n_3530);
  xnor g4595 (n_3501, n_1577, n_2447);
  or g4596 (n_3502, wc77, n_1577);
  not gc77 (wc77, n_2447);
  or g4597 (n_3504, wc78, n_1577);
  not gc78 (wc78, n_2448);
  and g4598 (n_3685, wc79, n_3538);
  not gc79 (wc79, n_3539);
  and g4599 (n_3679, n_3533, wc80);
  not gc80 (wc80, n_3541);
  not g4602 (Z[4], n_4101);
  or g4603 (n_4106, wc81, n_3541);
  not gc81 (wc81, n_3536);
  or g4604 (n_4109, wc82, n_3537);
  not gc82 (wc82, n_3538);
  and g4605 (n_3799, wc83, n_3536);
  not gc83 (wc83, n_3679);
  and g4606 (n_3686, n_3683, n_3533);
  xnor g4607 (Z[5], n_151, n_3530);
  or g4608 (n_4110, wc84, n_3547);
  not gc84 (wc84, n_3542);
  and g4609 (n_3688, wc85, n_3544);
  not gc85 (wc85, n_3545);
  and g4610 (n_3803, wc86, n_3685);
  not gc86 (wc86, n_3686);
  or g4611 (n_3884, wc87, n_3553);
  not gc87 (wc87, n_3691);
  or g4612 (n_4113, wc88, n_3543);
  not gc88 (wc88, n_3544);
  or g4613 (n_4115, wc89, n_3553);
  not gc89 (wc89, n_3548);
  and g4614 (n_3669, n_157, n_105);
  or g4615 (n_3670, n_157, n_105);
  and g4616 (n_3695, wc90, n_3550);
  not gc90 (wc90, n_3551);
  or g4619 (n_4118, wc91, n_3549);
  not gc91 (wc91, n_3550);
  and g4620 (n_3698, wc92, n_3556);
  not gc92 (wc92, n_3557);
  and g4621 (n_3886, wc93, n_3548);
  not gc93 (wc93, n_3689);
  and g4622 (n_3696, wc94, n_3693);
  not gc94 (wc94, n_3688);
  or g4623 (n_3882, n_3547, n_3803);
  or g4624 (n_3883, n_3803, wc95);
  not gc95 (wc95, n_3691);
  or g4625 (n_3887, n_3803, n_3884);
  xor g4626 (Z[7], n_4109, n_3799);
  xor g4627 (Z[8], n_4110, n_3803);
  or g4628 (n_4121, wc96, n_3559);
  not gc96 (wc96, n_3554);
  or g4629 (n_4124, wc97, n_3555);
  not gc97 (wc97, n_3556);
  or g4630 (n_4219, wc98, n_3671);
  not gc98 (wc98, n_3668);
  and g4631 (n_3705, wc99, n_3562);
  not gc99 (wc99, n_3563);
  and g4632 (n_3805, wc100, n_3695);
  not gc100 (wc100, n_3696);
  or g4633 (n_3812, wc101, n_3565);
  not gc101 (wc101, n_3701);
  and g4634 (n_3893, wc102, n_3701);
  not gc102 (wc102, n_3808);
  or g4635 (n_3889, n_3808, n_3803);
  or g4636 (n_3892, n_3803, wc103);
  not gc103 (wc103, n_3890);
  or g4637 (n_4126, wc104, n_3565);
  not gc104 (wc104, n_3560);
  or g4638 (n_4129, wc105, n_3561);
  not gc105 (wc105, n_3562);
  or g4639 (n_4130, wc106, n_3571);
  not gc106 (wc106, n_3566);
  or g4640 (n_4217, wc107, n_3663);
  not gc107 (wc107, n_3664);
  or g4641 (n_4222, wc108, n_3669);
  not gc108 (wc108, n_3670);
  and g4642 (n_3708, wc109, n_3568);
  not gc109 (wc109, n_3569);
  and g4643 (n_3788, wc110, n_3664);
  not gc110 (wc110, n_3665);
  and g4644 (n_3813, wc111, n_3560);
  not gc111 (wc111, n_3699);
  and g4645 (n_3706, wc112, n_3703);
  not gc112 (wc112, n_3698);
  or g4646 (n_4033, wc113, n_3671);
  not gc113 (wc113, n_3791);
  and g4647 (n_3810, wc114, n_3701);
  not gc114 (wc114, n_3805);
  or g4648 (n_3895, wc115, n_3803);
  not gc115 (wc115, n_3893);
  or g4649 (n_4133, wc116, n_3567);
  not gc116 (wc116, n_3568);
  or g4650 (n_4211, wc117, n_3657);
  not gc117 (wc117, n_3658);
  or g4651 (n_4214, wc118, n_3667);
  not gc118 (wc118, n_3662);
  and g4652 (n_3715, wc119, n_3574);
  not gc119 (wc119, n_3575);
  and g4653 (n_3718, wc120, n_3580);
  not gc120 (wc120, n_3581);
  and g4654 (n_3725, wc121, n_3586);
  not gc121 (wc121, n_3587);
  and g4655 (n_3778, wc122, n_3652);
  not gc122 (wc122, n_3653);
  and g4656 (n_3785, wc123, n_3658);
  not gc123 (wc123, n_3659);
  and g4657 (n_3817, wc124, n_3705);
  not gc124 (wc124, n_3706);
  or g4658 (n_3978, wc125, n_3577);
  not gc125 (wc125, n_3711);
  or g4659 (n_3827, wc126, n_3589);
  not gc126 (wc126, n_3721);
  or g4660 (n_3872, wc127, n_3661);
  not gc127 (wc127, n_3781);
  and g4661 (n_3891, wc128, n_3554);
  not gc128 (wc128, n_3806);
  and g4662 (n_3894, wc129, n_3698);
  not gc129 (wc129, n_3810);
  or g4663 (n_3898, n_3803, wc130);
  not gc130 (wc130, n_3896);
  or g4664 (n_3901, n_3803, wc131);
  not gc131 (wc131, n_3899);
  or g4665 (n_4135, wc132, n_3577);
  not gc132 (wc132, n_3572);
  or g4666 (n_4138, wc133, n_3573);
  not gc133 (wc133, n_3574);
  or g4667 (n_4141, wc134, n_3583);
  not gc134 (wc134, n_3578);
  or g4668 (n_4144, wc135, n_3579);
  not gc135 (wc135, n_3580);
  or g4669 (n_4146, wc136, n_3589);
  not gc136 (wc136, n_3584);
  or g4670 (n_4149, wc137, n_3585);
  not gc137 (wc137, n_3586);
  or g4671 (n_4203, wc138, n_3655);
  not gc138 (wc138, n_3650);
  or g4672 (n_4206, wc139, n_3651);
  not gc139 (wc139, n_3652);
  or g4673 (n_4208, wc140, n_3661);
  not gc140 (wc140, n_3656);
  and g4674 (n_3728, wc141, n_3592);
  not gc141 (wc141, n_3593);
  and g4675 (n_3775, wc142, n_3646);
  not gc142 (wc142, n_3647);
  and g4676 (n_3980, wc143, n_3572);
  not gc143 (wc143, n_3709);
  and g4677 (n_3716, wc144, n_3713);
  not gc144 (wc144, n_3708);
  and g4678 (n_3726, wc145, n_3723);
  not gc145 (wc145, n_3718);
  and g4679 (n_3786, wc146, n_3783);
  not gc146 (wc146, n_3778);
  and g4680 (n_4034, wc147, n_3668);
  not gc147 (wc147, n_3789);
  and g4681 (n_3897, n_3813, wc148);
  not gc148 (wc148, n_3814);
  and g4682 (n_3987, wc149, n_3721);
  not gc149 (wc149, n_3823);
  or g4683 (n_4151, wc150, n_3595);
  not gc150 (wc150, n_3590);
  or g4684 (n_4154, wc151, n_3591);
  not gc151 (wc151, n_3592);
  or g4685 (n_4197, wc152, n_3649);
  not gc152 (wc152, n_3644);
  or g4686 (n_4200, wc153, n_3645);
  not gc153 (wc153, n_3646);
  and g4687 (n_3735, wc154, n_3598);
  not gc154 (wc154, n_3599);
  and g4688 (n_3768, wc155, n_3640);
  not gc155 (wc155, n_3641);
  and g4689 (n_3820, wc156, n_3715);
  not gc156 (wc156, n_3716);
  and g4690 (n_3828, wc157, n_3584);
  not gc157 (wc157, n_3719);
  and g4691 (n_3832, wc158, n_3725);
  not gc158 (wc158, n_3726);
  or g4692 (n_3910, wc159, n_3601);
  not gc159 (wc159, n_3731);
  or g4693 (n_3946, wc160, n_3649);
  not gc160 (wc160, n_3771);
  and g4694 (n_3873, wc161, n_3656);
  not gc161 (wc161, n_3779);
  and g4695 (n_3877, wc162, n_3785);
  not gc162 (wc162, n_3786);
  and g4696 (n_3900, n_3817, wc163);
  not gc163 (wc163, n_3818);
  or g4697 (n_3994, wc164, n_3595);
  not gc164 (wc164, n_3905);
  or g4698 (n_4156, wc165, n_3601);
  not gc165 (wc165, n_3596);
  or g4699 (n_4159, wc166, n_3597);
  not gc166 (wc166, n_3598);
  or g4700 (n_4162, wc167, n_3607);
  not gc167 (wc167, n_3602);
  or g4701 (n_4167, wc168, n_3613);
  not gc168 (wc168, n_3608);
  or g4702 (n_4190, wc169, n_3633);
  not gc169 (wc169, n_3634);
  or g4703 (n_4192, wc170, n_3643);
  not gc170 (wc170, n_3638);
  or g4704 (n_4195, wc171, n_3639);
  not gc171 (wc171, n_3640);
  and g4705 (n_3738, wc172, n_3604);
  not gc172 (wc172, n_3605);
  and g4706 (n_3745, wc173, n_3610);
  not gc173 (wc173, n_3611);
  and g4707 (n_3748, wc174, n_3616);
  not gc174 (wc174, n_3617);
  and g4708 (n_3755, wc175, n_3622);
  not gc175 (wc175, n_3623);
  and g4709 (n_3758, wc176, n_3628);
  not gc176 (wc176, n_3629);
  and g4710 (n_3765, wc177, n_3634);
  not gc177 (wc177, n_3635);
  and g4711 (n_3911, wc178, n_3596);
  not gc178 (wc178, n_3729);
  and g4712 (n_3736, wc179, n_3733);
  not gc179 (wc179, n_3728);
  or g4713 (n_3842, wc180, n_3613);
  not gc180 (wc180, n_3741);
  or g4714 (n_4041, wc181, n_3625);
  not gc181 (wc181, n_3751);
  or g4715 (n_3857, wc182, n_3637);
  not gc182 (wc182, n_3761);
  and g4716 (n_3776, wc183, n_3773);
  not gc183 (wc183, n_3768);
  and g4717 (n_3825, wc184, n_3721);
  not gc184 (wc184, n_3820);
  and g4718 (n_3959, wc185, n_3781);
  not gc185 (wc185, n_3868);
  or g4719 (n_4165, wc186, n_3603);
  not gc186 (wc186, n_3604);
  or g4720 (n_4170, wc187, n_3609);
  not gc187 (wc187, n_3610);
  or g4721 (n_4171, wc188, n_3619);
  not gc188 (wc188, n_3614);
  or g4722 (n_4174, wc189, n_3615);
  not gc189 (wc189, n_3616);
  or g4723 (n_4176, wc190, n_3625);
  not gc190 (wc190, n_3620);
  or g4724 (n_4179, wc191, n_3621);
  not gc191 (wc191, n_3622);
  or g4725 (n_4182, wc192, n_3631);
  not gc192 (wc192, n_3626);
  or g4726 (n_4185, wc193, n_3627);
  not gc193 (wc193, n_3628);
  or g4727 (n_4187, wc194, n_3637);
  not gc194 (wc194, n_3632);
  and g4728 (n_3835, wc195, n_3735);
  not gc195 (wc195, n_3736);
  and g4729 (n_3746, wc196, n_3743);
  not gc196 (wc196, n_3738);
  and g4730 (n_3756, wc197, n_3753);
  not gc197 (wc197, n_3748);
  and g4731 (n_3766, wc198, n_3763);
  not gc198 (wc198, n_3758);
  and g4732 (n_3947, wc199, n_3644);
  not gc199 (wc199, n_3769);
  and g4733 (n_3865, wc200, n_3775);
  not gc200 (wc200, n_3776);
  and g4734 (n_3985, wc201, n_3578);
  not gc201 (wc201, n_3821);
  and g4735 (n_3988, wc202, n_3718);
  not gc202 (wc202, n_3825);
  and g4736 (n_3991, n_3828, wc203);
  not gc203 (wc203, n_3829);
  and g4737 (n_3902, n_3832, wc204);
  not gc204 (wc204, n_3833);
  and g4738 (n_3923, wc205, n_3741);
  not gc205 (wc205, n_3838);
  and g4739 (n_4050, wc206, n_3761);
  not gc206 (wc206, n_3853);
  or g4740 (n_4002, n_3910, wc207);
  not gc207 (wc207, n_3905);
  or g4741 (n_4006, wc208, n_3838);
  not gc208 (wc208, n_3905);
  or g4742 (n_3976, wc209, n_3571);
  not gc209 (wc209, n_3974);
  or g4743 (n_3981, n_3978, wc210);
  not gc210 (wc210, n_3974);
  or g4744 (n_3983, wc211, n_3823);
  not gc211 (wc211, n_3974);
  or g4745 (n_3997, n_3994, wc212);
  not gc212 (wc212, n_3974);
  or g4746 (n_4001, n_3998, wc213);
  not gc213 (wc213, n_3974);
  and g4747 (n_3843, wc214, n_3608);
  not gc214 (wc214, n_3739);
  and g4748 (n_3847, wc215, n_3745);
  not gc215 (wc215, n_3746);
  and g4749 (n_4043, wc216, n_3620);
  not gc216 (wc216, n_3749);
  and g4750 (n_3850, wc217, n_3755);
  not gc217 (wc217, n_3756);
  and g4751 (n_3858, wc218, n_3632);
  not gc218 (wc218, n_3759);
  and g4752 (n_3862, wc219, n_3765);
  not gc219 (wc219, n_3766);
  and g4753 (n_3840, wc220, n_3741);
  not gc220 (wc220, n_3835);
  and g4754 (n_3870, wc221, n_3781);
  not gc221 (wc221, n_3865);
  and g4755 (n_3908, wc222, n_3731);
  not gc222 (wc222, n_3902);
  and g4756 (n_3921, wc223, n_3918);
  not gc223 (wc223, n_3902);
  or g4757 (n_4057, wc224, n_3643);
  not gc224 (wc224, n_3941);
  or g4758 (n_4065, n_3946, wc225);
  not gc225 (wc225, n_3941);
  or g4759 (n_4069, wc226, n_3868);
  not gc226 (wc226, n_3941);
  and g4760 (n_3920, wc227, n_3602);
  not gc227 (wc227, n_3836);
  and g4761 (n_3925, wc228, n_3738);
  not gc228 (wc228, n_3840);
  and g4762 (n_3855, wc229, n_3761);
  not gc229 (wc229, n_3850);
  and g4763 (n_3956, wc230, n_3650);
  not gc230 (wc230, n_3866);
  and g4764 (n_3961, wc231, n_3778);
  not gc231 (wc231, n_3870);
  and g4765 (n_3966, n_3873, wc232);
  not gc232 (wc232, n_3874);
  and g4766 (n_3971, n_3877, wc233);
  not gc233 (wc233, n_3878);
  and g4767 (n_3996, wc234, n_3590);
  not gc234 (wc234, n_3903);
  and g4768 (n_4000, wc235, n_3728);
  not gc235 (wc235, n_3908);
  and g4769 (n_4004, n_3911, wc236);
  not gc236 (wc236, n_3912);
  and g4770 (n_4008, n_3835, wc237);
  not gc237 (wc237, n_3915);
  and g4771 (n_3926, n_3923, wc238);
  not gc238 (wc238, n_3902);
  and g4772 (n_3931, wc239, n_3928);
  not gc239 (wc239, n_3902);
  and g4773 (n_3936, wc240, n_3933);
  not gc240 (wc240, n_3902);
  or g4774 (n_4005, n_4002, wc241);
  not gc241 (wc241, n_3974);
  or g4775 (n_4009, n_4006, wc242);
  not gc242 (wc242, n_3974);
  or g4776 (n_4013, n_4010, wc243);
  not gc243 (wc243, n_3974);
  and g4777 (n_4090, wc244, n_3791);
  not gc244 (wc244, n_4029);
  and g4778 (n_3930, n_3843, wc245);
  not gc245 (wc245, n_3844);
  and g4779 (n_3935, n_3847, wc246);
  not gc246 (wc246, n_3848);
  and g4780 (n_4048, wc247, n_3626);
  not gc247 (wc247, n_3851);
  and g4781 (n_4051, wc248, n_3758);
  not gc248 (wc248, n_3855);
  and g4782 (n_4054, n_3858, wc249);
  not gc249 (wc249, n_3859);
  and g4783 (n_3938, n_3862, wc250);
  not gc250 (wc250, n_3863);
  or g4784 (n_4017, n_4014, wc251);
  not gc251 (wc251, n_3974);
  or g4785 (n_4021, n_4018, wc252);
  not gc252 (wc252, n_3974);
  or g4786 (n_4025, n_4022, wc253);
  not gc253 (wc253, n_3974);
  and g4787 (n_4012, n_3920, wc254);
  not gc254 (wc254, n_3921);
  and g4788 (n_4016, wc255, n_3925);
  not gc255 (wc255, n_3926);
  and g4789 (n_3944, wc256, n_3771);
  not gc256 (wc256, n_3938);
  and g4790 (n_3957, wc257, n_3954);
  not gc257 (wc257, n_3938);
  and g4791 (n_3962, wc258, n_3959);
  not gc258 (wc258, n_3938);
  and g4792 (n_3967, wc259, n_3964);
  not gc259 (wc259, n_3938);
  and g4793 (n_3972, wc260, n_3969);
  not gc260 (wc260, n_3938);
  and g4794 (n_4020, n_3930, wc261);
  not gc261 (wc261, n_3931);
  and g4795 (n_4024, n_3935, wc262);
  not gc262 (wc262, n_3936);
  and g4796 (n_4059, wc263, n_3638);
  not gc263 (wc263, n_3939);
  and g4797 (n_4063, wc264, n_3768);
  not gc264 (wc264, n_3944);
  and g4798 (n_4067, n_3947, wc265);
  not gc265 (wc265, n_3948);
  and g4799 (n_4071, n_3865, wc266);
  not gc266 (wc266, n_3951);
  and g4800 (n_4075, wc267, n_3956);
  not gc267 (wc267, n_3957);
  and g4801 (n_4079, wc268, n_3961);
  not gc268 (wc268, n_3962);
  and g4802 (n_4083, wc269, n_3966);
  not gc269 (wc269, n_3967);
  and g4803 (n_4026, wc270, n_3971);
  not gc270 (wc270, n_3972);
  and g4804 (n_4031, wc271, n_3791);
  not gc271 (wc271, n_4026);
  and g4805 (n_4088, wc272, n_3662);
  not gc272 (wc272, n_4027);
  and g4806 (n_4091, wc273, n_3788);
  not gc273 (wc273, n_4031);
  and g4807 (n_4094, n_4034, wc274);
  not gc274 (wc274, n_4035);
  or g4808 (n_4039, wc275, n_3619);
  not gc275 (wc275, n_4037);
  or g4809 (n_4044, n_4041, wc276);
  not gc276 (wc276, n_4037);
  or g4810 (n_4046, wc277, n_3853);
  not gc277 (wc277, n_4037);
  or g4811 (n_4060, n_4057, wc278);
  not gc278 (wc278, n_4037);
  or g4812 (n_4064, wc279, n_4061);
  not gc279 (wc279, n_4037);
  or g4813 (n_4068, n_4065, wc280);
  not gc280 (wc280, n_4037);
  or g4814 (n_4072, n_4069, wc281);
  not gc281 (wc281, n_4037);
  or g4815 (n_4076, wc282, n_4073);
  not gc282 (wc282, n_4037);
  or g4816 (n_4080, wc283, n_4077);
  not gc283 (wc283, n_4037);
  or g4817 (n_4084, wc284, n_4081);
  not gc284 (wc284, n_4037);
  or g4818 (n_4086, wc285, n_4029);
  not gc285 (wc285, n_4037);
endmodule

module mult_unsigned_GENERIC(A, B, Z);
  input [25:0] A, B;
  output [51:0] Z;
  wire [25:0] A, B;
  wire [51:0] Z;
  mult_unsigned_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

